magic
tech sky130A
magscale 1 2
timestamp 1636547095
<< viali >>
rect 1869 7497 1903 7531
rect 2513 7429 2547 7463
rect 5825 7429 5859 7463
rect 1961 7293 1995 7327
rect 4261 7293 4295 7327
rect 5181 7293 5215 7327
rect 6009 7293 6043 7327
rect 2697 7225 2731 7259
rect 4445 7157 4479 7191
rect 5365 7157 5399 7191
rect 2513 6817 2547 6851
rect 3157 6817 3191 6851
rect 4517 6817 4551 6851
rect 4261 6749 4295 6783
rect 2697 6681 2731 6715
rect 3341 6613 3375 6647
rect 5641 6613 5675 6647
rect 3157 6409 3191 6443
rect 2697 6341 2731 6375
rect 4537 6273 4571 6307
rect 5457 6273 5491 6307
rect 5549 6273 5583 6307
rect 1961 6205 1995 6239
rect 2513 6205 2547 6239
rect 1777 6137 1811 6171
rect 4270 6137 4304 6171
rect 4997 6069 5031 6103
rect 5365 6069 5399 6103
rect 3341 5865 3375 5899
rect 4261 5865 4295 5899
rect 2605 5729 2639 5763
rect 2789 5729 2823 5763
rect 3157 5729 3191 5763
rect 4445 5729 4479 5763
rect 4813 5729 4847 5763
rect 4997 5729 5031 5763
rect 5457 5729 5491 5763
rect 2881 5661 2915 5695
rect 2973 5661 3007 5695
rect 4629 5661 4663 5695
rect 4721 5661 4755 5695
rect 5549 5661 5583 5695
rect 1409 5321 1443 5355
rect 4721 5321 4755 5355
rect 5825 5321 5859 5355
rect 2789 5117 2823 5151
rect 5733 5117 5767 5151
rect 2544 5049 2578 5083
rect 3433 5049 3467 5083
rect 4261 4777 4295 4811
rect 5457 4777 5491 4811
rect 3249 4709 3283 4743
rect 5943 4709 5977 4743
rect 3157 4641 3191 4675
rect 4445 4641 4479 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 4997 4641 5031 4675
rect 5641 4641 5675 4675
rect 5733 4641 5767 4675
rect 5825 4641 5859 4675
rect 4721 4573 4755 4607
rect 6101 4573 6135 4607
rect 5181 4233 5215 4267
rect 3157 4097 3191 4131
rect 3249 4097 3283 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5733 4097 5767 4131
rect 2329 4029 2363 4063
rect 2973 4029 3007 4063
rect 3341 4029 3375 4063
rect 3525 4029 3559 4063
rect 5641 4029 5675 4063
rect 2145 3893 2179 3927
rect 2789 3893 2823 3927
rect 3985 3893 4019 3927
rect 4353 3893 4387 3927
rect 5549 3893 5583 3927
rect 4721 3689 4755 3723
rect 5181 3689 5215 3723
rect 3157 3621 3191 3655
rect 1777 3553 1811 3587
rect 2605 3553 2639 3587
rect 5089 3553 5123 3587
rect 6101 3553 6135 3587
rect 5365 3485 5399 3519
rect 1961 3417 1995 3451
rect 2421 3349 2455 3383
rect 3249 3349 3283 3383
rect 5917 3349 5951 3383
rect 3709 3145 3743 3179
rect 4261 3145 4295 3179
rect 5457 3077 5491 3111
rect 2329 3009 2363 3043
rect 4905 3009 4939 3043
rect 1685 2941 1719 2975
rect 2596 2941 2630 2975
rect 4454 2941 4488 2975
rect 4747 2941 4781 2975
rect 5457 2941 5491 2975
rect 5733 2941 5767 2975
rect 4537 2873 4571 2907
rect 4629 2873 4663 2907
rect 1869 2805 1903 2839
rect 4261 2601 4295 2635
rect 5365 2601 5399 2635
rect 2329 2533 2363 2567
rect 3157 2533 3191 2567
rect 3341 2533 3375 2567
rect 4629 2533 4663 2567
rect 4747 2533 4781 2567
rect 5733 2533 5767 2567
rect 1593 2465 1627 2499
rect 2973 2465 3007 2499
rect 4445 2465 4479 2499
rect 4537 2465 4571 2499
rect 4905 2465 4939 2499
rect 5549 2465 5583 2499
rect 5641 2465 5675 2499
rect 5851 2465 5885 2499
rect 6009 2465 6043 2499
rect 1777 2329 1811 2363
rect 2421 2261 2455 2295
<< metal1 >>
rect 1104 7642 6808 7664
rect 1104 7590 1932 7642
rect 1984 7590 1996 7642
rect 2048 7590 2060 7642
rect 2112 7590 2124 7642
rect 2176 7590 3834 7642
rect 3886 7590 3898 7642
rect 3950 7590 3962 7642
rect 4014 7590 4026 7642
rect 4078 7590 5735 7642
rect 5787 7590 5799 7642
rect 5851 7590 5863 7642
rect 5915 7590 5927 7642
rect 5979 7590 6808 7642
rect 1104 7568 6808 7590
rect 1857 7531 1915 7537
rect 1857 7497 1869 7531
rect 1903 7528 1915 7531
rect 2774 7528 2780 7540
rect 1903 7500 2780 7528
rect 1903 7497 1915 7500
rect 1857 7491 1915 7497
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 2501 7463 2559 7469
rect 2501 7460 2513 7463
rect 1820 7432 2513 7460
rect 1820 7420 1826 7432
rect 2501 7429 2513 7432
rect 2547 7429 2559 7463
rect 2501 7423 2559 7429
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 5813 7463 5871 7469
rect 5813 7460 5825 7463
rect 5408 7432 5825 7460
rect 5408 7420 5414 7432
rect 5813 7429 5825 7432
rect 5859 7429 5871 7463
rect 5813 7423 5871 7429
rect 7374 7392 7380 7404
rect 5184 7364 7380 7392
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7324 2007 7327
rect 2774 7324 2780 7336
rect 1995 7296 2780 7324
rect 1995 7293 2007 7296
rect 1949 7287 2007 7293
rect 2774 7284 2780 7296
rect 2832 7284 2838 7336
rect 3694 7284 3700 7336
rect 3752 7324 3758 7336
rect 5184 7333 5212 7364
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 4249 7327 4307 7333
rect 4249 7324 4261 7327
rect 3752 7296 4261 7324
rect 3752 7284 3758 7296
rect 4249 7293 4261 7296
rect 4295 7293 4307 7327
rect 4249 7287 4307 7293
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 5442 7284 5448 7336
rect 5500 7324 5506 7336
rect 5997 7327 6055 7333
rect 5997 7324 6009 7327
rect 5500 7296 6009 7324
rect 5500 7284 5506 7296
rect 5997 7293 6009 7296
rect 6043 7293 6055 7327
rect 5997 7287 6055 7293
rect 2685 7259 2743 7265
rect 2685 7225 2697 7259
rect 2731 7256 2743 7259
rect 3234 7256 3240 7268
rect 2731 7228 3240 7256
rect 2731 7225 2743 7228
rect 2685 7219 2743 7225
rect 3234 7216 3240 7228
rect 3292 7216 3298 7268
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 5626 7188 5632 7200
rect 5399 7160 5632 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 1104 7098 6808 7120
rect 1104 7046 2883 7098
rect 2935 7046 2947 7098
rect 2999 7046 3011 7098
rect 3063 7046 3075 7098
rect 3127 7046 4784 7098
rect 4836 7046 4848 7098
rect 4900 7046 4912 7098
rect 4964 7046 4976 7098
rect 5028 7046 6808 7098
rect 1104 7024 6808 7046
rect 3252 6888 4660 6916
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 3145 6851 3203 6857
rect 3145 6817 3157 6851
rect 3191 6848 3203 6851
rect 3252 6848 3280 6888
rect 3191 6820 3280 6848
rect 3191 6817 3203 6820
rect 3145 6811 3203 6817
rect 3326 6808 3332 6860
rect 3384 6848 3390 6860
rect 4505 6851 4563 6857
rect 4505 6848 4517 6851
rect 3384 6820 4517 6848
rect 3384 6808 3390 6820
rect 4505 6817 4517 6820
rect 4551 6817 4563 6851
rect 4632 6848 4660 6888
rect 5534 6848 5540 6860
rect 4632 6820 5540 6848
rect 4505 6811 4563 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 2685 6715 2743 6721
rect 2685 6681 2697 6715
rect 2731 6712 2743 6715
rect 4264 6712 4292 6743
rect 2731 6684 4292 6712
rect 2731 6681 2743 6684
rect 2685 6675 2743 6681
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 4154 6644 4160 6656
rect 3375 6616 4160 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4264 6644 4292 6684
rect 4522 6644 4528 6656
rect 4264 6616 4528 6644
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5316 6616 5641 6644
rect 5316 6604 5322 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 1104 6554 6808 6576
rect 1104 6502 1932 6554
rect 1984 6502 1996 6554
rect 2048 6502 2060 6554
rect 2112 6502 2124 6554
rect 2176 6502 3834 6554
rect 3886 6502 3898 6554
rect 3950 6502 3962 6554
rect 4014 6502 4026 6554
rect 4078 6502 5735 6554
rect 5787 6502 5799 6554
rect 5851 6502 5863 6554
rect 5915 6502 5927 6554
rect 5979 6502 6808 6554
rect 1104 6480 6808 6502
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3234 6440 3240 6452
rect 3191 6412 3240 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 5074 6440 5080 6452
rect 4396 6412 5080 6440
rect 4396 6400 4402 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 2685 6375 2743 6381
rect 2685 6341 2697 6375
rect 2731 6372 2743 6375
rect 3510 6372 3516 6384
rect 2731 6344 3516 6372
rect 2731 6341 2743 6344
rect 2685 6335 2743 6341
rect 3510 6332 3516 6344
rect 3568 6332 3574 6384
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5445 6307 5503 6313
rect 5445 6304 5457 6307
rect 5408 6276 5457 6304
rect 5408 6264 5414 6276
rect 5445 6273 5457 6276
rect 5491 6273 5503 6307
rect 5445 6267 5503 6273
rect 5534 6264 5540 6316
rect 5592 6304 5598 6316
rect 5592 6276 5637 6304
rect 5592 6264 5598 6276
rect 1394 6196 1400 6248
rect 1452 6236 1458 6248
rect 1949 6239 2007 6245
rect 1949 6236 1961 6239
rect 1452 6208 1961 6236
rect 1452 6196 1458 6208
rect 1949 6205 1961 6208
rect 1995 6205 2007 6239
rect 1949 6199 2007 6205
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 1762 6168 1768 6180
rect 1723 6140 1768 6168
rect 1762 6128 1768 6140
rect 1820 6128 1826 6180
rect 2516 6168 2544 6199
rect 2774 6196 2780 6248
rect 2832 6236 2838 6248
rect 5258 6236 5264 6248
rect 2832 6208 5264 6236
rect 2832 6196 2838 6208
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 3602 6168 3608 6180
rect 2516 6140 3608 6168
rect 3602 6128 3608 6140
rect 3660 6128 3666 6180
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 4258 6171 4316 6177
rect 4258 6168 4270 6171
rect 4212 6140 4270 6168
rect 4212 6128 4218 6140
rect 4258 6137 4270 6140
rect 4304 6137 4316 6171
rect 4258 6131 4316 6137
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 4985 6103 5043 6109
rect 4985 6100 4997 6103
rect 4580 6072 4997 6100
rect 4580 6060 4586 6072
rect 4985 6069 4997 6072
rect 5031 6069 5043 6103
rect 5350 6100 5356 6112
rect 5311 6072 5356 6100
rect 4985 6063 5043 6069
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 1104 6010 6808 6032
rect 1104 5958 2883 6010
rect 2935 5958 2947 6010
rect 2999 5958 3011 6010
rect 3063 5958 3075 6010
rect 3127 5958 4784 6010
rect 4836 5958 4848 6010
rect 4900 5958 4912 6010
rect 4964 5958 4976 6010
rect 5028 5958 6808 6010
rect 1104 5936 6808 5958
rect 3326 5896 3332 5908
rect 3287 5868 3332 5896
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 4249 5899 4307 5905
rect 4249 5896 4261 5899
rect 4212 5868 4261 5896
rect 4212 5856 4218 5868
rect 4249 5865 4261 5868
rect 4295 5865 4307 5899
rect 4522 5896 4528 5908
rect 4249 5859 4307 5865
rect 4448 5868 4528 5896
rect 4448 5828 4476 5868
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 4264 5800 4476 5828
rect 2593 5763 2651 5769
rect 2593 5729 2605 5763
rect 2639 5729 2651 5763
rect 2593 5723 2651 5729
rect 2608 5624 2636 5723
rect 2774 5720 2780 5772
rect 2832 5760 2838 5772
rect 3145 5763 3203 5769
rect 2832 5732 2877 5760
rect 2832 5720 2838 5732
rect 3145 5729 3157 5763
rect 3191 5760 3203 5763
rect 4264 5760 4292 5800
rect 5074 5788 5080 5840
rect 5132 5828 5138 5840
rect 5132 5800 5488 5828
rect 5132 5788 5138 5800
rect 3191 5732 4292 5760
rect 3191 5729 3203 5732
rect 3145 5723 3203 5729
rect 4338 5720 4344 5772
rect 4396 5760 4402 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 4396 5732 4445 5760
rect 4396 5720 4402 5732
rect 4433 5729 4445 5732
rect 4479 5729 4491 5763
rect 4798 5760 4804 5772
rect 4759 5732 4804 5760
rect 4433 5723 4491 5729
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5760 5043 5763
rect 5166 5760 5172 5772
rect 5031 5732 5172 5760
rect 5031 5729 5043 5732
rect 4985 5723 5043 5729
rect 5166 5720 5172 5732
rect 5224 5720 5230 5772
rect 5460 5769 5488 5800
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 2866 5692 2872 5704
rect 2827 5664 2872 5692
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 4614 5692 4620 5704
rect 3007 5664 4620 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 5184 5692 5212 5720
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5184 5664 5549 5692
rect 4709 5655 4767 5661
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 4154 5624 4160 5636
rect 2608 5596 4160 5624
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 4724 5624 4752 5655
rect 4632 5596 4752 5624
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 4632 5556 4660 5596
rect 2924 5528 4660 5556
rect 2924 5516 2930 5528
rect 1104 5466 6808 5488
rect 1104 5414 1932 5466
rect 1984 5414 1996 5466
rect 2048 5414 2060 5466
rect 2112 5414 2124 5466
rect 2176 5414 3834 5466
rect 3886 5414 3898 5466
rect 3950 5414 3962 5466
rect 4014 5414 4026 5466
rect 4078 5414 5735 5466
rect 5787 5414 5799 5466
rect 5851 5414 5863 5466
rect 5915 5414 5927 5466
rect 5979 5414 6808 5466
rect 1104 5392 6808 5414
rect 1394 5352 1400 5364
rect 1355 5324 1400 5352
rect 1394 5312 1400 5324
rect 1452 5312 1458 5364
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 4709 5355 4767 5361
rect 4709 5352 4721 5355
rect 2556 5324 4721 5352
rect 2556 5312 2562 5324
rect 4709 5321 4721 5324
rect 4755 5321 4767 5355
rect 4709 5315 4767 5321
rect 5534 5312 5540 5364
rect 5592 5352 5598 5364
rect 5813 5355 5871 5361
rect 5813 5352 5825 5355
rect 5592 5324 5825 5352
rect 5592 5312 5598 5324
rect 5813 5321 5825 5324
rect 5859 5321 5871 5355
rect 5813 5315 5871 5321
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 5721 5151 5779 5157
rect 2832 5120 2877 5148
rect 2832 5108 2838 5120
rect 5721 5117 5733 5151
rect 5767 5148 5779 5151
rect 5810 5148 5816 5160
rect 5767 5120 5816 5148
rect 5767 5117 5779 5120
rect 5721 5111 5779 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 2532 5083 2590 5089
rect 2532 5049 2544 5083
rect 2578 5080 2590 5083
rect 3326 5080 3332 5092
rect 2578 5052 3332 5080
rect 2578 5049 2590 5052
rect 2532 5043 2590 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 3418 5040 3424 5092
rect 3476 5080 3482 5092
rect 3476 5052 3521 5080
rect 3476 5040 3482 5052
rect 1104 4922 6808 4944
rect 1104 4870 2883 4922
rect 2935 4870 2947 4922
rect 2999 4870 3011 4922
rect 3063 4870 3075 4922
rect 3127 4870 4784 4922
rect 4836 4870 4848 4922
rect 4900 4870 4912 4922
rect 4964 4870 4976 4922
rect 5028 4870 6808 4922
rect 1104 4848 6808 4870
rect 3326 4768 3332 4820
rect 3384 4808 3390 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 3384 4780 4261 4808
rect 3384 4768 3390 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 5408 4780 5457 4808
rect 5408 4768 5414 4780
rect 5445 4777 5457 4780
rect 5491 4777 5503 4811
rect 5445 4771 5503 4777
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 3237 4743 3295 4749
rect 3237 4740 3249 4743
rect 3108 4712 3249 4740
rect 3108 4700 3114 4712
rect 3237 4709 3249 4712
rect 3283 4740 3295 4743
rect 5074 4740 5080 4752
rect 3283 4712 4660 4740
rect 3283 4709 3295 4712
rect 3237 4703 3295 4709
rect 4632 4684 4660 4712
rect 4816 4712 5080 4740
rect 3145 4675 3203 4681
rect 3145 4641 3157 4675
rect 3191 4672 3203 4675
rect 4433 4675 4491 4681
rect 3191 4644 3280 4672
rect 3191 4641 3203 4644
rect 3145 4635 3203 4641
rect 3252 4616 3280 4644
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4522 4672 4528 4684
rect 4479 4644 4528 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 4614 4632 4620 4684
rect 4672 4672 4678 4684
rect 4816 4681 4844 4712
rect 5074 4700 5080 4712
rect 5132 4740 5138 4752
rect 5931 4743 5989 4749
rect 5931 4740 5943 4743
rect 5132 4712 5943 4740
rect 5132 4700 5138 4712
rect 5931 4709 5943 4712
rect 5977 4709 5989 4743
rect 5931 4703 5989 4709
rect 4801 4675 4859 4681
rect 4672 4644 4717 4672
rect 4672 4632 4678 4644
rect 4801 4641 4813 4675
rect 4847 4641 4859 4675
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4801 4635 4859 4641
rect 4908 4644 4997 4672
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 4709 4607 4767 4613
rect 4709 4604 4721 4607
rect 3292 4576 4721 4604
rect 3292 4564 3298 4576
rect 4709 4573 4721 4576
rect 4755 4573 4767 4607
rect 4709 4567 4767 4573
rect 1394 4496 1400 4548
rect 1452 4536 1458 4548
rect 4816 4536 4844 4635
rect 1452 4508 4844 4536
rect 1452 4496 1458 4508
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4908 4468 4936 4644
rect 4985 4641 4997 4644
rect 5031 4672 5043 4675
rect 5166 4672 5172 4684
rect 5031 4644 5172 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5626 4672 5632 4684
rect 5587 4644 5632 4672
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 5721 4675 5779 4681
rect 5721 4641 5733 4675
rect 5767 4641 5779 4675
rect 5721 4635 5779 4641
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 5736 4604 5764 4635
rect 5810 4632 5816 4684
rect 5868 4672 5874 4684
rect 6270 4672 6276 4684
rect 5868 4644 6276 4672
rect 5868 4632 5874 4644
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 5500 4576 5764 4604
rect 6089 4607 6147 4613
rect 5500 4564 5506 4576
rect 6089 4573 6101 4607
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 5626 4496 5632 4548
rect 5684 4536 5690 4548
rect 6104 4536 6132 4567
rect 5684 4508 6132 4536
rect 5684 4496 5690 4508
rect 4212 4440 4936 4468
rect 4212 4428 4218 4440
rect 1104 4378 6808 4400
rect 1104 4326 1932 4378
rect 1984 4326 1996 4378
rect 2048 4326 2060 4378
rect 2112 4326 2124 4378
rect 2176 4326 3834 4378
rect 3886 4326 3898 4378
rect 3950 4326 3962 4378
rect 4014 4326 4026 4378
rect 4078 4326 5735 4378
rect 5787 4326 5799 4378
rect 5851 4326 5863 4378
rect 5915 4326 5927 4378
rect 5979 4326 6808 4378
rect 1104 4304 6808 4326
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 5169 4267 5227 4273
rect 5169 4264 5181 4267
rect 4580 4236 5181 4264
rect 4580 4224 4586 4236
rect 5169 4233 5181 4236
rect 5215 4233 5227 4267
rect 5169 4227 5227 4233
rect 3050 4088 3056 4140
rect 3108 4128 3114 4140
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 3108 4100 3157 4128
rect 3108 4088 3114 4100
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3234 4088 3240 4140
rect 3292 4128 3298 4140
rect 3292 4100 3337 4128
rect 3292 4088 3298 4100
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4304 4100 4445 4128
rect 4304 4088 4310 4100
rect 4433 4097 4445 4100
rect 4479 4128 4491 4131
rect 4522 4128 4528 4140
rect 4479 4100 4528 4128
rect 4479 4097 4491 4100
rect 4433 4091 4491 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 5534 4128 5540 4140
rect 4663 4100 5540 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 5534 4088 5540 4100
rect 5592 4128 5598 4140
rect 5721 4131 5779 4137
rect 5721 4128 5733 4131
rect 5592 4100 5733 4128
rect 5592 4088 5598 4100
rect 5721 4097 5733 4100
rect 5767 4097 5779 4131
rect 5721 4091 5779 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2498 4060 2504 4072
rect 2363 4032 2504 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2774 4060 2780 4072
rect 2746 4020 2780 4060
rect 2832 4020 2838 4072
rect 2961 4063 3019 4069
rect 2961 4029 2973 4063
rect 3007 4029 3019 4063
rect 3326 4060 3332 4072
rect 3287 4032 3332 4060
rect 2961 4023 3019 4029
rect 2746 3992 2774 4020
rect 2148 3964 2774 3992
rect 2148 3933 2176 3964
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 2648 3896 2789 3924
rect 2648 3884 2654 3896
rect 2777 3893 2789 3896
rect 2823 3893 2835 3927
rect 2976 3924 3004 4023
rect 3326 4020 3332 4032
rect 3384 4020 3390 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 4154 4060 4160 4072
rect 3559 4032 4160 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 4154 4020 4160 4032
rect 4212 4020 4218 4072
rect 5258 4020 5264 4072
rect 5316 4060 5322 4072
rect 5629 4063 5687 4069
rect 5629 4060 5641 4063
rect 5316 4032 5641 4060
rect 5316 4020 5322 4032
rect 5629 4029 5641 4032
rect 5675 4029 5687 4063
rect 5629 4023 5687 4029
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 2976 3896 3985 3924
rect 2777 3887 2835 3893
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 4246 3884 4252 3936
rect 4304 3924 4310 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4304 3896 4353 3924
rect 4304 3884 4310 3896
rect 4341 3893 4353 3896
rect 4387 3893 4399 3927
rect 4341 3887 4399 3893
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 5224 3896 5549 3924
rect 5224 3884 5230 3896
rect 5537 3893 5549 3896
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 1104 3834 6808 3856
rect 1104 3782 2883 3834
rect 2935 3782 2947 3834
rect 2999 3782 3011 3834
rect 3063 3782 3075 3834
rect 3127 3782 4784 3834
rect 4836 3782 4848 3834
rect 4900 3782 4912 3834
rect 4964 3782 4976 3834
rect 5028 3782 6808 3834
rect 1104 3760 6808 3782
rect 4338 3680 4344 3732
rect 4396 3720 4402 3732
rect 4709 3723 4767 3729
rect 4709 3720 4721 3723
rect 4396 3692 4721 3720
rect 4396 3680 4402 3692
rect 4709 3689 4721 3692
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 5132 3692 5181 3720
rect 5132 3680 5138 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 3145 3655 3203 3661
rect 3145 3621 3157 3655
rect 3191 3652 3203 3655
rect 3510 3652 3516 3664
rect 3191 3624 3516 3652
rect 3191 3621 3203 3624
rect 3145 3615 3203 3621
rect 3510 3612 3516 3624
rect 3568 3612 3574 3664
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2593 3587 2651 3593
rect 2593 3553 2605 3587
rect 2639 3553 2651 3587
rect 5074 3584 5080 3596
rect 5035 3556 5080 3584
rect 2593 3547 2651 3553
rect 2608 3516 2636 3547
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 6086 3584 6092 3596
rect 6047 3556 6092 3584
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 4154 3516 4160 3528
rect 2608 3488 4160 3516
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5534 3516 5540 3528
rect 5399 3488 5540 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5534 3476 5540 3488
rect 5592 3516 5598 3528
rect 6178 3516 6184 3528
rect 5592 3488 6184 3516
rect 5592 3476 5598 3488
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 4522 3448 4528 3460
rect 1995 3420 4528 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 4522 3408 4528 3420
rect 4580 3408 4586 3460
rect 2406 3380 2412 3392
rect 2367 3352 2412 3380
rect 2406 3340 2412 3352
rect 2464 3340 2470 3392
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 4614 3380 4620 3392
rect 3283 3352 4620 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5592 3352 5917 3380
rect 5592 3340 5598 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 5905 3343 5963 3349
rect 1104 3290 6808 3312
rect 1104 3238 1932 3290
rect 1984 3238 1996 3290
rect 2048 3238 2060 3290
rect 2112 3238 2124 3290
rect 2176 3238 3834 3290
rect 3886 3238 3898 3290
rect 3950 3238 3962 3290
rect 4014 3238 4026 3290
rect 4078 3238 5735 3290
rect 5787 3238 5799 3290
rect 5851 3238 5863 3290
rect 5915 3238 5927 3290
rect 5979 3238 6808 3290
rect 1104 3216 6808 3238
rect 2682 3176 2688 3188
rect 2332 3148 2688 3176
rect 2332 3049 2360 3148
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3694 3176 3700 3188
rect 3384 3148 3700 3176
rect 3384 3136 3390 3148
rect 3694 3136 3700 3148
rect 3752 3136 3758 3188
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 4430 3068 4436 3120
rect 4488 3068 4494 3120
rect 5445 3111 5503 3117
rect 5445 3108 5457 3111
rect 4908 3080 5457 3108
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 474 2932 480 2984
rect 532 2972 538 2984
rect 2590 2981 2596 2984
rect 1673 2975 1731 2981
rect 1673 2972 1685 2975
rect 532 2944 1685 2972
rect 532 2932 538 2944
rect 1673 2941 1685 2944
rect 1719 2941 1731 2975
rect 2584 2972 2596 2981
rect 2551 2944 2596 2972
rect 1673 2935 1731 2941
rect 2584 2935 2596 2944
rect 2590 2932 2596 2935
rect 2648 2932 2654 2984
rect 4448 2981 4476 3068
rect 4522 3000 4528 3052
rect 4580 3000 4586 3052
rect 4908 3049 4936 3080
rect 5445 3077 5457 3080
rect 5491 3108 5503 3111
rect 5626 3108 5632 3120
rect 5491 3080 5632 3108
rect 5491 3077 5503 3080
rect 5445 3071 5503 3077
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 5718 3068 5724 3120
rect 5776 3108 5782 3120
rect 6270 3108 6276 3120
rect 5776 3080 6276 3108
rect 5776 3068 5782 3080
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 4442 2975 4500 2981
rect 4442 2941 4454 2975
rect 4488 2941 4500 2975
rect 4540 2972 4568 3000
rect 4735 2975 4793 2981
rect 4735 2972 4747 2975
rect 4540 2944 4747 2972
rect 4442 2935 4500 2941
rect 4735 2941 4747 2944
rect 4781 2941 4793 2975
rect 5442 2972 5448 2984
rect 5403 2944 5448 2972
rect 4735 2935 4793 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5721 2975 5779 2981
rect 5721 2941 5733 2975
rect 5767 2972 5779 2975
rect 6178 2972 6184 2984
rect 5767 2944 6184 2972
rect 5767 2941 5779 2944
rect 5721 2935 5779 2941
rect 6178 2932 6184 2944
rect 6236 2932 6242 2984
rect 4338 2904 4344 2916
rect 1872 2876 4344 2904
rect 1872 2845 1900 2876
rect 4338 2864 4344 2876
rect 4396 2864 4402 2916
rect 4522 2904 4528 2916
rect 4483 2876 4528 2904
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2904 4675 2907
rect 4890 2904 4896 2916
rect 4663 2876 4896 2904
rect 4663 2873 4675 2876
rect 4617 2867 4675 2873
rect 4890 2864 4896 2876
rect 4948 2904 4954 2916
rect 4948 2876 5764 2904
rect 4948 2864 4954 2876
rect 5736 2848 5764 2876
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2805 1915 2839
rect 1857 2799 1915 2805
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 3326 2836 3332 2848
rect 2372 2808 3332 2836
rect 2372 2796 2378 2808
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 5166 2836 5172 2848
rect 4304 2808 5172 2836
rect 4304 2796 4310 2808
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 5718 2796 5724 2848
rect 5776 2796 5782 2848
rect 1104 2746 6808 2768
rect 1104 2694 2883 2746
rect 2935 2694 2947 2746
rect 2999 2694 3011 2746
rect 3063 2694 3075 2746
rect 3127 2694 4784 2746
rect 4836 2694 4848 2746
rect 4900 2694 4912 2746
rect 4964 2694 4976 2746
rect 5028 2694 6808 2746
rect 1104 2672 6808 2694
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4430 2592 4436 2644
rect 4488 2592 4494 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5132 2604 5365 2632
rect 5132 2592 5138 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5626 2632 5632 2644
rect 5539 2604 5632 2632
rect 5353 2595 5411 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2406 2564 2412 2576
rect 2363 2536 2412 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2406 2524 2412 2536
rect 2464 2564 2470 2576
rect 3145 2567 3203 2573
rect 3145 2564 3157 2567
rect 2464 2536 3157 2564
rect 2464 2524 2470 2536
rect 3145 2533 3157 2536
rect 3191 2533 3203 2567
rect 3145 2527 3203 2533
rect 3234 2524 3240 2576
rect 3292 2564 3298 2576
rect 3329 2567 3387 2573
rect 3329 2564 3341 2567
rect 3292 2536 3341 2564
rect 3292 2524 3298 2536
rect 3329 2533 3341 2536
rect 3375 2533 3387 2567
rect 4448 2564 4476 2592
rect 4617 2567 4675 2573
rect 4617 2564 4629 2567
rect 3329 2527 3387 2533
rect 3988 2536 4629 2564
rect 1581 2499 1639 2505
rect 1581 2465 1593 2499
rect 1627 2465 1639 2499
rect 1581 2459 1639 2465
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2496 3019 2499
rect 3418 2496 3424 2508
rect 3007 2468 3424 2496
rect 3007 2465 3019 2468
rect 2961 2459 3019 2465
rect 1596 2428 1624 2459
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3786 2428 3792 2440
rect 1596 2400 3792 2428
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 1765 2363 1823 2369
rect 1765 2329 1777 2363
rect 1811 2360 1823 2363
rect 3694 2360 3700 2372
rect 1811 2332 3700 2360
rect 1811 2329 1823 2332
rect 1765 2323 1823 2329
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 2409 2295 2467 2301
rect 2409 2261 2421 2295
rect 2455 2292 2467 2295
rect 3988 2292 4016 2536
rect 4617 2533 4629 2536
rect 4663 2533 4675 2567
rect 4617 2527 4675 2533
rect 4706 2524 4712 2576
rect 4764 2573 4770 2576
rect 4764 2567 4793 2573
rect 4781 2533 4793 2567
rect 5552 2564 5580 2604
rect 5626 2592 5632 2604
rect 5684 2632 5690 2644
rect 5684 2604 6040 2632
rect 5684 2592 5690 2604
rect 5718 2564 5724 2576
rect 4764 2527 4793 2533
rect 4908 2536 5580 2564
rect 5679 2536 5724 2564
rect 4764 2524 4770 2527
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4396 2468 4445 2496
rect 4396 2456 4402 2468
rect 4433 2465 4445 2468
rect 4479 2465 4491 2499
rect 4433 2459 4491 2465
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 4908 2505 4936 2536
rect 5718 2524 5724 2536
rect 5776 2524 5782 2576
rect 4893 2499 4951 2505
rect 4580 2468 4673 2496
rect 4580 2456 4586 2468
rect 4893 2465 4905 2499
rect 4939 2465 4951 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 4893 2459 4951 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6012 2505 6040 2604
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5839 2499 5897 2505
rect 5839 2496 5851 2499
rect 5629 2459 5687 2465
rect 5736 2468 5851 2496
rect 4540 2428 4568 2456
rect 4540 2400 4660 2428
rect 4062 2320 4068 2372
rect 4120 2320 4126 2372
rect 4632 2360 4660 2400
rect 5442 2388 5448 2440
rect 5500 2428 5506 2440
rect 5644 2428 5672 2459
rect 5500 2400 5672 2428
rect 5500 2388 5506 2400
rect 5460 2360 5488 2388
rect 4632 2332 5488 2360
rect 2455 2264 4016 2292
rect 4080 2292 4108 2320
rect 5736 2292 5764 2468
rect 5839 2465 5851 2468
rect 5885 2465 5897 2499
rect 5839 2459 5897 2465
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 4080 2264 5764 2292
rect 2455 2261 2467 2264
rect 2409 2255 2467 2261
rect 1104 2202 6808 2224
rect 1104 2150 1932 2202
rect 1984 2150 1996 2202
rect 2048 2150 2060 2202
rect 2112 2150 2124 2202
rect 2176 2150 3834 2202
rect 3886 2150 3898 2202
rect 3950 2150 3962 2202
rect 4014 2150 4026 2202
rect 4078 2150 5735 2202
rect 5787 2150 5799 2202
rect 5851 2150 5863 2202
rect 5915 2150 5927 2202
rect 5979 2150 6808 2202
rect 1104 2128 6808 2150
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 5994 1272 6000 1284
rect 3660 1244 6000 1272
rect 3660 1232 3666 1244
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
<< via1 >>
rect 1932 7590 1984 7642
rect 1996 7590 2048 7642
rect 2060 7590 2112 7642
rect 2124 7590 2176 7642
rect 3834 7590 3886 7642
rect 3898 7590 3950 7642
rect 3962 7590 4014 7642
rect 4026 7590 4078 7642
rect 5735 7590 5787 7642
rect 5799 7590 5851 7642
rect 5863 7590 5915 7642
rect 5927 7590 5979 7642
rect 2780 7488 2832 7540
rect 1768 7420 1820 7472
rect 5356 7420 5408 7472
rect 2780 7284 2832 7336
rect 3700 7284 3752 7336
rect 7380 7352 7432 7404
rect 5448 7284 5500 7336
rect 3240 7216 3292 7268
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 5632 7148 5684 7200
rect 2883 7046 2935 7098
rect 2947 7046 2999 7098
rect 3011 7046 3063 7098
rect 3075 7046 3127 7098
rect 4784 7046 4836 7098
rect 4848 7046 4900 7098
rect 4912 7046 4964 7098
rect 4976 7046 5028 7098
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 3332 6808 3384 6860
rect 5540 6808 5592 6860
rect 4160 6604 4212 6656
rect 4528 6604 4580 6656
rect 5264 6604 5316 6656
rect 1932 6502 1984 6554
rect 1996 6502 2048 6554
rect 2060 6502 2112 6554
rect 2124 6502 2176 6554
rect 3834 6502 3886 6554
rect 3898 6502 3950 6554
rect 3962 6502 4014 6554
rect 4026 6502 4078 6554
rect 5735 6502 5787 6554
rect 5799 6502 5851 6554
rect 5863 6502 5915 6554
rect 5927 6502 5979 6554
rect 3240 6400 3292 6452
rect 4344 6400 4396 6452
rect 5080 6400 5132 6452
rect 3516 6332 3568 6384
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5356 6264 5408 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 1400 6196 1452 6248
rect 1768 6171 1820 6180
rect 1768 6137 1777 6171
rect 1777 6137 1811 6171
rect 1811 6137 1820 6171
rect 1768 6128 1820 6137
rect 2780 6196 2832 6248
rect 5264 6196 5316 6248
rect 3608 6128 3660 6180
rect 4160 6128 4212 6180
rect 4528 6060 4580 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 2883 5958 2935 6010
rect 2947 5958 2999 6010
rect 3011 5958 3063 6010
rect 3075 5958 3127 6010
rect 4784 5958 4836 6010
rect 4848 5958 4900 6010
rect 4912 5958 4964 6010
rect 4976 5958 5028 6010
rect 3332 5899 3384 5908
rect 3332 5865 3341 5899
rect 3341 5865 3375 5899
rect 3375 5865 3384 5899
rect 3332 5856 3384 5865
rect 4160 5856 4212 5908
rect 4528 5856 4580 5908
rect 2780 5763 2832 5772
rect 2780 5729 2789 5763
rect 2789 5729 2823 5763
rect 2823 5729 2832 5763
rect 2780 5720 2832 5729
rect 5080 5788 5132 5840
rect 4344 5720 4396 5772
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 5172 5720 5224 5772
rect 2872 5695 2924 5704
rect 2872 5661 2881 5695
rect 2881 5661 2915 5695
rect 2915 5661 2924 5695
rect 2872 5652 2924 5661
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4160 5584 4212 5636
rect 2872 5516 2924 5568
rect 1932 5414 1984 5466
rect 1996 5414 2048 5466
rect 2060 5414 2112 5466
rect 2124 5414 2176 5466
rect 3834 5414 3886 5466
rect 3898 5414 3950 5466
rect 3962 5414 4014 5466
rect 4026 5414 4078 5466
rect 5735 5414 5787 5466
rect 5799 5414 5851 5466
rect 5863 5414 5915 5466
rect 5927 5414 5979 5466
rect 1400 5355 1452 5364
rect 1400 5321 1409 5355
rect 1409 5321 1443 5355
rect 1443 5321 1452 5355
rect 1400 5312 1452 5321
rect 2504 5312 2556 5364
rect 5540 5312 5592 5364
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 5816 5108 5868 5160
rect 3332 5040 3384 5092
rect 3424 5083 3476 5092
rect 3424 5049 3433 5083
rect 3433 5049 3467 5083
rect 3467 5049 3476 5083
rect 3424 5040 3476 5049
rect 2883 4870 2935 4922
rect 2947 4870 2999 4922
rect 3011 4870 3063 4922
rect 3075 4870 3127 4922
rect 4784 4870 4836 4922
rect 4848 4870 4900 4922
rect 4912 4870 4964 4922
rect 4976 4870 5028 4922
rect 3332 4768 3384 4820
rect 5356 4768 5408 4820
rect 3056 4700 3108 4752
rect 4528 4632 4580 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 5080 4700 5132 4752
rect 4620 4632 4672 4641
rect 3240 4564 3292 4616
rect 1400 4496 1452 4548
rect 4160 4428 4212 4480
rect 5172 4632 5224 4684
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 5448 4564 5500 4616
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6276 4632 6328 4684
rect 5632 4496 5684 4548
rect 1932 4326 1984 4378
rect 1996 4326 2048 4378
rect 2060 4326 2112 4378
rect 2124 4326 2176 4378
rect 3834 4326 3886 4378
rect 3898 4326 3950 4378
rect 3962 4326 4014 4378
rect 4026 4326 4078 4378
rect 5735 4326 5787 4378
rect 5799 4326 5851 4378
rect 5863 4326 5915 4378
rect 5927 4326 5979 4378
rect 4528 4224 4580 4276
rect 3056 4088 3108 4140
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 4252 4088 4304 4140
rect 4528 4088 4580 4140
rect 5540 4088 5592 4140
rect 2504 4020 2556 4072
rect 2780 4020 2832 4072
rect 3332 4063 3384 4072
rect 2596 3884 2648 3936
rect 3332 4029 3341 4063
rect 3341 4029 3375 4063
rect 3375 4029 3384 4063
rect 3332 4020 3384 4029
rect 4160 4020 4212 4072
rect 5264 4020 5316 4072
rect 4252 3884 4304 3936
rect 5172 3884 5224 3936
rect 2883 3782 2935 3834
rect 2947 3782 2999 3834
rect 3011 3782 3063 3834
rect 3075 3782 3127 3834
rect 4784 3782 4836 3834
rect 4848 3782 4900 3834
rect 4912 3782 4964 3834
rect 4976 3782 5028 3834
rect 4344 3680 4396 3732
rect 5080 3680 5132 3732
rect 3516 3612 3568 3664
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 4160 3476 4212 3528
rect 5540 3476 5592 3528
rect 6184 3476 6236 3528
rect 4528 3408 4580 3460
rect 2412 3383 2464 3392
rect 2412 3349 2421 3383
rect 2421 3349 2455 3383
rect 2455 3349 2464 3383
rect 2412 3340 2464 3349
rect 4620 3340 4672 3392
rect 5540 3340 5592 3392
rect 1932 3238 1984 3290
rect 1996 3238 2048 3290
rect 2060 3238 2112 3290
rect 2124 3238 2176 3290
rect 3834 3238 3886 3290
rect 3898 3238 3950 3290
rect 3962 3238 4014 3290
rect 4026 3238 4078 3290
rect 5735 3238 5787 3290
rect 5799 3238 5851 3290
rect 5863 3238 5915 3290
rect 5927 3238 5979 3290
rect 2688 3136 2740 3188
rect 3332 3136 3384 3188
rect 3700 3179 3752 3188
rect 3700 3145 3709 3179
rect 3709 3145 3743 3179
rect 3743 3145 3752 3179
rect 3700 3136 3752 3145
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 4436 3068 4488 3120
rect 480 2932 532 2984
rect 2596 2975 2648 2984
rect 2596 2941 2630 2975
rect 2630 2941 2648 2975
rect 2596 2932 2648 2941
rect 4528 3000 4580 3052
rect 5632 3068 5684 3120
rect 5724 3068 5776 3120
rect 6276 3068 6328 3120
rect 5448 2975 5500 2984
rect 5448 2941 5457 2975
rect 5457 2941 5491 2975
rect 5491 2941 5500 2975
rect 5448 2932 5500 2941
rect 6184 2932 6236 2984
rect 4344 2864 4396 2916
rect 4528 2907 4580 2916
rect 4528 2873 4537 2907
rect 4537 2873 4571 2907
rect 4571 2873 4580 2907
rect 4528 2864 4580 2873
rect 4896 2864 4948 2916
rect 2320 2796 2372 2848
rect 3332 2796 3384 2848
rect 4252 2796 4304 2848
rect 5172 2796 5224 2848
rect 5724 2796 5776 2848
rect 2883 2694 2935 2746
rect 2947 2694 2999 2746
rect 3011 2694 3063 2746
rect 3075 2694 3127 2746
rect 4784 2694 4836 2746
rect 4848 2694 4900 2746
rect 4912 2694 4964 2746
rect 4976 2694 5028 2746
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 4436 2592 4488 2644
rect 5080 2592 5132 2644
rect 2412 2524 2464 2576
rect 3240 2524 3292 2576
rect 3424 2456 3476 2508
rect 3792 2388 3844 2440
rect 3700 2320 3752 2372
rect 4712 2567 4764 2576
rect 4712 2533 4747 2567
rect 4747 2533 4764 2567
rect 5632 2592 5684 2644
rect 5724 2567 5776 2576
rect 4712 2524 4764 2533
rect 4344 2456 4396 2508
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 5724 2533 5733 2567
rect 5733 2533 5767 2567
rect 5767 2533 5776 2567
rect 5724 2524 5776 2533
rect 4528 2456 4580 2465
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 4068 2320 4120 2372
rect 5448 2388 5500 2440
rect 1932 2150 1984 2202
rect 1996 2150 2048 2202
rect 2060 2150 2112 2202
rect 2124 2150 2176 2202
rect 3834 2150 3886 2202
rect 3898 2150 3950 2202
rect 3962 2150 4014 2202
rect 4026 2150 4078 2202
rect 5735 2150 5787 2202
rect 5799 2150 5851 2202
rect 5863 2150 5915 2202
rect 5927 2150 5979 2202
rect 3608 1232 3660 1284
rect 6000 1232 6052 1284
<< metal2 >>
rect 1858 9343 1914 10143
rect 3698 9343 3754 10143
rect 5538 9343 5594 10143
rect 7378 9343 7434 10143
rect 1872 7834 1900 9343
rect 2778 8936 2834 8945
rect 2778 8871 2834 8880
rect 1780 7806 1900 7834
rect 1780 7478 1808 7806
rect 1906 7644 2202 7664
rect 1962 7642 1986 7644
rect 2042 7642 2066 7644
rect 2122 7642 2146 7644
rect 1984 7590 1986 7642
rect 2048 7590 2060 7642
rect 2122 7590 2124 7642
rect 1962 7588 1986 7590
rect 2042 7588 2066 7590
rect 2122 7588 2146 7590
rect 1906 7568 2202 7588
rect 2792 7546 2820 8871
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 3712 7342 3740 9343
rect 3808 7644 4104 7664
rect 3864 7642 3888 7644
rect 3944 7642 3968 7644
rect 4024 7642 4048 7644
rect 3886 7590 3888 7642
rect 3950 7590 3962 7642
rect 4024 7590 4026 7642
rect 3864 7588 3888 7590
rect 3944 7588 3968 7590
rect 4024 7588 4048 7590
rect 3808 7568 4104 7588
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 1906 6556 2202 6576
rect 1962 6554 1986 6556
rect 2042 6554 2066 6556
rect 2122 6554 2146 6556
rect 1984 6502 1986 6554
rect 2048 6502 2060 6554
rect 2122 6502 2124 6554
rect 1962 6500 1986 6502
rect 2042 6500 2066 6502
rect 2122 6500 2146 6502
rect 1906 6480 2202 6500
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1766 6216 1822 6225
rect 1412 5370 1440 6190
rect 1766 6151 1768 6160
rect 1820 6151 1822 6160
rect 1768 6122 1820 6128
rect 1906 5468 2202 5488
rect 1962 5466 1986 5468
rect 2042 5466 2066 5468
rect 2122 5466 2146 5468
rect 1984 5414 1986 5466
rect 2048 5414 2060 5466
rect 2122 5414 2124 5466
rect 1962 5412 1986 5414
rect 2042 5412 2066 5414
rect 2122 5412 2146 5414
rect 1906 5392 2202 5412
rect 2516 5370 2544 6802
rect 2792 6254 2820 7278
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 2857 7100 3153 7120
rect 2913 7098 2937 7100
rect 2993 7098 3017 7100
rect 3073 7098 3097 7100
rect 2935 7046 2937 7098
rect 2999 7046 3011 7098
rect 3073 7046 3075 7098
rect 2913 7044 2937 7046
rect 2993 7044 3017 7046
rect 3073 7044 3097 7046
rect 2857 7024 3153 7044
rect 3252 6458 3280 7210
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 2780 6248 2832 6254
rect 2780 6190 2832 6196
rect 2792 5778 2820 6190
rect 2857 6012 3153 6032
rect 2913 6010 2937 6012
rect 2993 6010 3017 6012
rect 3073 6010 3097 6012
rect 2935 5958 2937 6010
rect 2999 5958 3011 6010
rect 3073 5958 3075 6010
rect 2913 5956 2937 5958
rect 2993 5956 3017 5958
rect 3073 5956 3097 5958
rect 2857 5936 3153 5956
rect 3252 5817 3280 6394
rect 3344 5914 3372 6802
rect 4160 6656 4212 6662
rect 4212 6604 4384 6610
rect 4160 6598 4384 6604
rect 4172 6582 4384 6598
rect 3808 6556 4104 6576
rect 3864 6554 3888 6556
rect 3944 6554 3968 6556
rect 4024 6554 4048 6556
rect 3886 6502 3888 6554
rect 3950 6502 3962 6554
rect 4024 6502 4026 6554
rect 3864 6500 3888 6502
rect 3944 6500 3968 6502
rect 4024 6500 4048 6502
rect 3808 6480 4104 6500
rect 4356 6458 4384 6582
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3238 5808 3294 5817
rect 2780 5772 2832 5778
rect 3238 5743 3294 5752
rect 2780 5714 2832 5720
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5574 2912 5646
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 1412 4554 1440 5306
rect 1400 4548 1452 4554
rect 1400 4490 1452 4496
rect 1906 4380 2202 4400
rect 1962 4378 1986 4380
rect 2042 4378 2066 4380
rect 2122 4378 2146 4380
rect 1984 4326 1986 4378
rect 2048 4326 2060 4378
rect 2122 4326 2124 4378
rect 1962 4324 1986 4326
rect 2042 4324 2066 4326
rect 2122 4324 2146 4326
rect 1906 4304 2202 4324
rect 2516 4078 2544 5306
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2884 5114 2912 5510
rect 2792 4078 2820 5102
rect 2884 5086 3280 5114
rect 2857 4924 3153 4944
rect 2913 4922 2937 4924
rect 2993 4922 3017 4924
rect 3073 4922 3097 4924
rect 2935 4870 2937 4922
rect 2999 4870 3011 4922
rect 3073 4870 3075 4922
rect 2913 4868 2937 4870
rect 2993 4868 3017 4870
rect 3073 4868 3097 4870
rect 2857 4848 3153 4868
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3068 4146 3096 4694
rect 3252 4622 3280 5086
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3344 4826 3372 5034
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4146 3280 4558
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3505 1808 3538
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 2412 3392 2464 3398
rect 2412 3334 2464 3340
rect 1906 3292 2202 3312
rect 1962 3290 1986 3292
rect 2042 3290 2066 3292
rect 2122 3290 2146 3292
rect 1984 3238 1986 3290
rect 2048 3238 2060 3290
rect 2122 3238 2124 3290
rect 1962 3236 1986 3238
rect 2042 3236 2066 3238
rect 2122 3236 2146 3238
rect 1906 3216 2202 3236
rect 480 2984 532 2990
rect 480 2926 532 2932
rect 492 800 520 2926
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 1906 2204 2202 2224
rect 1962 2202 1986 2204
rect 2042 2202 2066 2204
rect 2122 2202 2146 2204
rect 1984 2150 1986 2202
rect 2048 2150 2060 2202
rect 2122 2150 2124 2202
rect 1962 2148 1986 2150
rect 2042 2148 2066 2150
rect 2122 2148 2146 2150
rect 1906 2128 2202 2148
rect 2332 800 2360 2790
rect 2424 2582 2452 3334
rect 2608 2990 2636 3878
rect 2792 3210 2820 4014
rect 2857 3836 3153 3856
rect 2913 3834 2937 3836
rect 2993 3834 3017 3836
rect 3073 3834 3097 3836
rect 2935 3782 2937 3834
rect 2999 3782 3011 3834
rect 3073 3782 3075 3834
rect 2913 3780 2937 3782
rect 2993 3780 3017 3782
rect 3073 3780 3097 3782
rect 2857 3760 3153 3780
rect 2700 3194 2820 3210
rect 2688 3188 2820 3194
rect 2740 3182 2820 3188
rect 2688 3130 2740 3136
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2857 2748 3153 2768
rect 2913 2746 2937 2748
rect 2993 2746 3017 2748
rect 3073 2746 3097 2748
rect 2935 2694 2937 2746
rect 2999 2694 3011 2746
rect 3073 2694 3075 2746
rect 2913 2692 2937 2694
rect 2993 2692 3017 2694
rect 3073 2692 3097 2694
rect 2857 2672 3153 2692
rect 3252 2582 3280 4082
rect 3332 4072 3384 4078
rect 3332 4014 3384 4020
rect 3344 3194 3372 4014
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3332 2848 3384 2854
rect 3436 2836 3464 5034
rect 3528 3670 3556 6326
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 3384 2808 3464 2836
rect 3332 2790 3384 2796
rect 3528 2774 3556 3606
rect 3436 2746 3556 2774
rect 2412 2576 2464 2582
rect 2412 2518 2464 2524
rect 3240 2576 3292 2582
rect 3240 2518 3292 2524
rect 3436 2514 3464 2746
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3620 1290 3648 6122
rect 4172 5914 4200 6122
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4250 5808 4306 5817
rect 4250 5743 4306 5752
rect 4344 5772 4396 5778
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 3808 5468 4104 5488
rect 3864 5466 3888 5468
rect 3944 5466 3968 5468
rect 4024 5466 4048 5468
rect 3886 5414 3888 5466
rect 3950 5414 3962 5466
rect 4024 5414 4026 5466
rect 3864 5412 3888 5414
rect 3944 5412 3968 5414
rect 4024 5412 4048 5414
rect 3808 5392 4104 5412
rect 4172 4486 4200 5578
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3808 4380 4104 4400
rect 3864 4378 3888 4380
rect 3944 4378 3968 4380
rect 4024 4378 4048 4380
rect 3886 4326 3888 4378
rect 3950 4326 3962 4378
rect 4024 4326 4026 4378
rect 3864 4324 3888 4326
rect 3944 4324 3968 4326
rect 4024 4324 4048 4326
rect 3808 4304 4104 4324
rect 4172 4078 4200 4422
rect 4264 4146 4292 5743
rect 4344 5714 4396 5720
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 4072 4212 4078
rect 4160 4014 4212 4020
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 3808 3292 4104 3312
rect 3864 3290 3888 3292
rect 3944 3290 3968 3292
rect 4024 3290 4048 3292
rect 3886 3238 3888 3290
rect 3950 3238 3962 3290
rect 4024 3238 4026 3290
rect 3864 3236 3888 3238
rect 3944 3236 3968 3238
rect 4024 3236 4048 3238
rect 3808 3216 4104 3236
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3712 2564 3740 3130
rect 3712 2536 4108 2564
rect 3804 2446 3832 2536
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4080 2378 4108 2536
rect 3700 2372 3752 2378
rect 3700 2314 3752 2320
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 478 0 534 800
rect 2318 0 2374 800
rect 3712 785 3740 2314
rect 3808 2204 4104 2224
rect 3864 2202 3888 2204
rect 3944 2202 3968 2204
rect 4024 2202 4048 2204
rect 3886 2150 3888 2202
rect 3950 2150 3962 2202
rect 4024 2150 4026 2202
rect 3864 2148 3888 2150
rect 3944 2148 3968 2150
rect 4024 2148 4048 2150
rect 3808 2128 4104 2148
rect 4172 800 4200 3470
rect 4264 3194 4292 3878
rect 4356 3738 4384 5714
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4448 3126 4476 7142
rect 4758 7100 5054 7120
rect 4814 7098 4838 7100
rect 4894 7098 4918 7100
rect 4974 7098 4998 7100
rect 4836 7046 4838 7098
rect 4900 7046 4912 7098
rect 4974 7046 4976 7098
rect 4814 7044 4838 7046
rect 4894 7044 4918 7046
rect 4974 7044 4998 7046
rect 4758 7024 5054 7044
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4540 6322 4568 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5914 4568 6054
rect 4758 6012 5054 6032
rect 4814 6010 4838 6012
rect 4894 6010 4918 6012
rect 4974 6010 4998 6012
rect 4836 5958 4838 6010
rect 4900 5958 4912 6010
rect 4974 5958 4976 6010
rect 4814 5956 4838 5958
rect 4894 5956 4918 5958
rect 4974 5956 4998 5958
rect 4758 5936 5054 5956
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 5092 5846 5120 6394
rect 5276 6254 5304 6598
rect 5368 6322 5396 7414
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5264 6248 5316 6254
rect 5460 6225 5488 7278
rect 5552 6866 5580 9343
rect 5709 7644 6005 7664
rect 5765 7642 5789 7644
rect 5845 7642 5869 7644
rect 5925 7642 5949 7644
rect 5787 7590 5789 7642
rect 5851 7590 5863 7642
rect 5925 7590 5927 7642
rect 5765 7588 5789 7590
rect 5845 7588 5869 7590
rect 5925 7588 5949 7590
rect 5709 7568 6005 7588
rect 7392 7410 7420 9343
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5540 6316 5592 6322
rect 5540 6258 5592 6264
rect 5264 6190 5316 6196
rect 5446 6216 5502 6225
rect 5080 5840 5132 5846
rect 4802 5808 4858 5817
rect 5080 5782 5132 5788
rect 4802 5743 4804 5752
rect 4856 5743 4858 5752
rect 5172 5772 5224 5778
rect 4804 5714 4856 5720
rect 5172 5714 5224 5720
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4632 4690 4660 5646
rect 4758 4924 5054 4944
rect 4814 4922 4838 4924
rect 4894 4922 4918 4924
rect 4974 4922 4998 4924
rect 4836 4870 4838 4922
rect 4900 4870 4912 4922
rect 4974 4870 4976 4922
rect 4814 4868 4838 4870
rect 4894 4868 4918 4870
rect 4974 4868 4998 4870
rect 4758 4848 5054 4868
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 4620 4684 4672 4690
rect 4620 4626 4672 4632
rect 4540 4282 4568 4626
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4528 4140 4580 4146
rect 4580 4100 4660 4128
rect 4528 4082 4580 4088
rect 4632 3482 4660 4100
rect 4758 3836 5054 3856
rect 4814 3834 4838 3836
rect 4894 3834 4918 3836
rect 4974 3834 4998 3836
rect 4836 3782 4838 3834
rect 4900 3782 4912 3834
rect 4974 3782 4976 3834
rect 4814 3780 4838 3782
rect 4894 3780 4918 3782
rect 4974 3780 4998 3782
rect 4758 3760 5054 3780
rect 5092 3738 5120 4694
rect 5184 4690 5212 5714
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5276 4078 5304 6190
rect 5446 6151 5502 6160
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 4826 5396 6054
rect 5552 5370 5580 6258
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4528 3460 4580 3466
rect 4632 3454 4752 3482
rect 4528 3402 4580 3408
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4540 3058 4568 3402
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4528 3052 4580 3058
rect 4528 2994 4580 3000
rect 4632 2938 4660 3334
rect 4540 2922 4660 2938
rect 4344 2916 4396 2922
rect 4344 2858 4396 2864
rect 4528 2916 4660 2922
rect 4580 2910 4660 2916
rect 4528 2858 4580 2864
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4264 2650 4292 2790
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4356 2514 4384 2858
rect 4434 2816 4490 2825
rect 4434 2751 4490 2760
rect 4448 2650 4476 2751
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4540 2514 4568 2858
rect 4724 2836 4752 3454
rect 4894 2952 4950 2961
rect 4894 2887 4896 2896
rect 4948 2887 4950 2896
rect 4896 2858 4948 2864
rect 4632 2808 4752 2836
rect 4632 2564 4660 2808
rect 4758 2748 5054 2768
rect 4814 2746 4838 2748
rect 4894 2746 4918 2748
rect 4974 2746 4998 2748
rect 4836 2694 4838 2746
rect 4900 2694 4912 2746
rect 4974 2694 4976 2746
rect 4814 2692 4838 2694
rect 4894 2692 4918 2694
rect 4974 2692 4998 2694
rect 4758 2672 5054 2692
rect 5092 2650 5120 3538
rect 5184 2854 5212 3878
rect 5460 2990 5488 4558
rect 5552 4146 5580 5306
rect 5644 4690 5672 7142
rect 5709 6556 6005 6576
rect 5765 6554 5789 6556
rect 5845 6554 5869 6556
rect 5925 6554 5949 6556
rect 5787 6502 5789 6554
rect 5851 6502 5863 6554
rect 5925 6502 5927 6554
rect 5765 6500 5789 6502
rect 5845 6500 5869 6502
rect 5925 6500 5949 6502
rect 5709 6480 6005 6500
rect 5709 5468 6005 5488
rect 5765 5466 5789 5468
rect 5845 5466 5869 5468
rect 5925 5466 5949 5468
rect 5787 5414 5789 5466
rect 5851 5414 5863 5466
rect 5925 5414 5927 5466
rect 5765 5412 5789 5414
rect 5845 5412 5869 5414
rect 5925 5412 5949 5414
rect 5709 5392 6005 5412
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4690 5856 5102
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 5632 4548 5684 4554
rect 5632 4490 5684 4496
rect 5540 4140 5592 4146
rect 5540 4082 5592 4088
rect 5552 3534 5580 4082
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 4712 2576 4764 2582
rect 4632 2536 4712 2564
rect 4712 2518 4764 2524
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 5460 2446 5488 2926
rect 5552 2514 5580 3334
rect 5644 3126 5672 4490
rect 5709 4380 6005 4400
rect 5765 4378 5789 4380
rect 5845 4378 5869 4380
rect 5925 4378 5949 4380
rect 5787 4326 5789 4378
rect 5851 4326 5863 4378
rect 5925 4326 5927 4378
rect 5765 4324 5789 4326
rect 5845 4324 5869 4326
rect 5925 4324 5949 4326
rect 5709 4304 6005 4324
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6104 3505 6132 3538
rect 6184 3528 6236 3534
rect 6090 3496 6146 3505
rect 6184 3470 6236 3476
rect 6090 3431 6146 3440
rect 5709 3292 6005 3312
rect 5765 3290 5789 3292
rect 5845 3290 5869 3292
rect 5925 3290 5949 3292
rect 5787 3238 5789 3290
rect 5851 3238 5863 3290
rect 5925 3238 5927 3290
rect 5765 3236 5789 3238
rect 5845 3236 5869 3238
rect 5925 3236 5949 3238
rect 5709 3216 6005 3236
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5644 2650 5672 3062
rect 5736 2854 5764 3062
rect 6196 2990 6224 3470
rect 6288 3126 6316 4626
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6184 2984 6236 2990
rect 6184 2926 6236 2932
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5736 2582 5764 2790
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5709 2204 6005 2224
rect 5765 2202 5789 2204
rect 5845 2202 5869 2204
rect 5925 2202 5949 2204
rect 5787 2150 5789 2202
rect 5851 2150 5863 2202
rect 5925 2150 5927 2202
rect 5765 2148 5789 2150
rect 5845 2148 5869 2150
rect 5925 2148 5949 2150
rect 5709 2128 6005 2148
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 6012 800 6040 1226
rect 3698 776 3754 785
rect 3698 711 3754 720
rect 4158 0 4214 800
rect 5998 0 6054 800
<< via2 >>
rect 2778 8880 2834 8936
rect 1906 7642 1962 7644
rect 1986 7642 2042 7644
rect 2066 7642 2122 7644
rect 2146 7642 2202 7644
rect 1906 7590 1932 7642
rect 1932 7590 1962 7642
rect 1986 7590 1996 7642
rect 1996 7590 2042 7642
rect 2066 7590 2112 7642
rect 2112 7590 2122 7642
rect 2146 7590 2176 7642
rect 2176 7590 2202 7642
rect 1906 7588 1962 7590
rect 1986 7588 2042 7590
rect 2066 7588 2122 7590
rect 2146 7588 2202 7590
rect 3808 7642 3864 7644
rect 3888 7642 3944 7644
rect 3968 7642 4024 7644
rect 4048 7642 4104 7644
rect 3808 7590 3834 7642
rect 3834 7590 3864 7642
rect 3888 7590 3898 7642
rect 3898 7590 3944 7642
rect 3968 7590 4014 7642
rect 4014 7590 4024 7642
rect 4048 7590 4078 7642
rect 4078 7590 4104 7642
rect 3808 7588 3864 7590
rect 3888 7588 3944 7590
rect 3968 7588 4024 7590
rect 4048 7588 4104 7590
rect 1906 6554 1962 6556
rect 1986 6554 2042 6556
rect 2066 6554 2122 6556
rect 2146 6554 2202 6556
rect 1906 6502 1932 6554
rect 1932 6502 1962 6554
rect 1986 6502 1996 6554
rect 1996 6502 2042 6554
rect 2066 6502 2112 6554
rect 2112 6502 2122 6554
rect 2146 6502 2176 6554
rect 2176 6502 2202 6554
rect 1906 6500 1962 6502
rect 1986 6500 2042 6502
rect 2066 6500 2122 6502
rect 2146 6500 2202 6502
rect 1766 6180 1822 6216
rect 1766 6160 1768 6180
rect 1768 6160 1820 6180
rect 1820 6160 1822 6180
rect 1906 5466 1962 5468
rect 1986 5466 2042 5468
rect 2066 5466 2122 5468
rect 2146 5466 2202 5468
rect 1906 5414 1932 5466
rect 1932 5414 1962 5466
rect 1986 5414 1996 5466
rect 1996 5414 2042 5466
rect 2066 5414 2112 5466
rect 2112 5414 2122 5466
rect 2146 5414 2176 5466
rect 2176 5414 2202 5466
rect 1906 5412 1962 5414
rect 1986 5412 2042 5414
rect 2066 5412 2122 5414
rect 2146 5412 2202 5414
rect 2857 7098 2913 7100
rect 2937 7098 2993 7100
rect 3017 7098 3073 7100
rect 3097 7098 3153 7100
rect 2857 7046 2883 7098
rect 2883 7046 2913 7098
rect 2937 7046 2947 7098
rect 2947 7046 2993 7098
rect 3017 7046 3063 7098
rect 3063 7046 3073 7098
rect 3097 7046 3127 7098
rect 3127 7046 3153 7098
rect 2857 7044 2913 7046
rect 2937 7044 2993 7046
rect 3017 7044 3073 7046
rect 3097 7044 3153 7046
rect 2857 6010 2913 6012
rect 2937 6010 2993 6012
rect 3017 6010 3073 6012
rect 3097 6010 3153 6012
rect 2857 5958 2883 6010
rect 2883 5958 2913 6010
rect 2937 5958 2947 6010
rect 2947 5958 2993 6010
rect 3017 5958 3063 6010
rect 3063 5958 3073 6010
rect 3097 5958 3127 6010
rect 3127 5958 3153 6010
rect 2857 5956 2913 5958
rect 2937 5956 2993 5958
rect 3017 5956 3073 5958
rect 3097 5956 3153 5958
rect 3808 6554 3864 6556
rect 3888 6554 3944 6556
rect 3968 6554 4024 6556
rect 4048 6554 4104 6556
rect 3808 6502 3834 6554
rect 3834 6502 3864 6554
rect 3888 6502 3898 6554
rect 3898 6502 3944 6554
rect 3968 6502 4014 6554
rect 4014 6502 4024 6554
rect 4048 6502 4078 6554
rect 4078 6502 4104 6554
rect 3808 6500 3864 6502
rect 3888 6500 3944 6502
rect 3968 6500 4024 6502
rect 4048 6500 4104 6502
rect 3238 5752 3294 5808
rect 1906 4378 1962 4380
rect 1986 4378 2042 4380
rect 2066 4378 2122 4380
rect 2146 4378 2202 4380
rect 1906 4326 1932 4378
rect 1932 4326 1962 4378
rect 1986 4326 1996 4378
rect 1996 4326 2042 4378
rect 2066 4326 2112 4378
rect 2112 4326 2122 4378
rect 2146 4326 2176 4378
rect 2176 4326 2202 4378
rect 1906 4324 1962 4326
rect 1986 4324 2042 4326
rect 2066 4324 2122 4326
rect 2146 4324 2202 4326
rect 2857 4922 2913 4924
rect 2937 4922 2993 4924
rect 3017 4922 3073 4924
rect 3097 4922 3153 4924
rect 2857 4870 2883 4922
rect 2883 4870 2913 4922
rect 2937 4870 2947 4922
rect 2947 4870 2993 4922
rect 3017 4870 3063 4922
rect 3063 4870 3073 4922
rect 3097 4870 3127 4922
rect 3127 4870 3153 4922
rect 2857 4868 2913 4870
rect 2937 4868 2993 4870
rect 3017 4868 3073 4870
rect 3097 4868 3153 4870
rect 1766 3440 1822 3496
rect 1906 3290 1962 3292
rect 1986 3290 2042 3292
rect 2066 3290 2122 3292
rect 2146 3290 2202 3292
rect 1906 3238 1932 3290
rect 1932 3238 1962 3290
rect 1986 3238 1996 3290
rect 1996 3238 2042 3290
rect 2066 3238 2112 3290
rect 2112 3238 2122 3290
rect 2146 3238 2176 3290
rect 2176 3238 2202 3290
rect 1906 3236 1962 3238
rect 1986 3236 2042 3238
rect 2066 3236 2122 3238
rect 2146 3236 2202 3238
rect 1906 2202 1962 2204
rect 1986 2202 2042 2204
rect 2066 2202 2122 2204
rect 2146 2202 2202 2204
rect 1906 2150 1932 2202
rect 1932 2150 1962 2202
rect 1986 2150 1996 2202
rect 1996 2150 2042 2202
rect 2066 2150 2112 2202
rect 2112 2150 2122 2202
rect 2146 2150 2176 2202
rect 2176 2150 2202 2202
rect 1906 2148 1962 2150
rect 1986 2148 2042 2150
rect 2066 2148 2122 2150
rect 2146 2148 2202 2150
rect 2857 3834 2913 3836
rect 2937 3834 2993 3836
rect 3017 3834 3073 3836
rect 3097 3834 3153 3836
rect 2857 3782 2883 3834
rect 2883 3782 2913 3834
rect 2937 3782 2947 3834
rect 2947 3782 2993 3834
rect 3017 3782 3063 3834
rect 3063 3782 3073 3834
rect 3097 3782 3127 3834
rect 3127 3782 3153 3834
rect 2857 3780 2913 3782
rect 2937 3780 2993 3782
rect 3017 3780 3073 3782
rect 3097 3780 3153 3782
rect 2857 2746 2913 2748
rect 2937 2746 2993 2748
rect 3017 2746 3073 2748
rect 3097 2746 3153 2748
rect 2857 2694 2883 2746
rect 2883 2694 2913 2746
rect 2937 2694 2947 2746
rect 2947 2694 2993 2746
rect 3017 2694 3063 2746
rect 3063 2694 3073 2746
rect 3097 2694 3127 2746
rect 3127 2694 3153 2746
rect 2857 2692 2913 2694
rect 2937 2692 2993 2694
rect 3017 2692 3073 2694
rect 3097 2692 3153 2694
rect 4250 5752 4306 5808
rect 3808 5466 3864 5468
rect 3888 5466 3944 5468
rect 3968 5466 4024 5468
rect 4048 5466 4104 5468
rect 3808 5414 3834 5466
rect 3834 5414 3864 5466
rect 3888 5414 3898 5466
rect 3898 5414 3944 5466
rect 3968 5414 4014 5466
rect 4014 5414 4024 5466
rect 4048 5414 4078 5466
rect 4078 5414 4104 5466
rect 3808 5412 3864 5414
rect 3888 5412 3944 5414
rect 3968 5412 4024 5414
rect 4048 5412 4104 5414
rect 3808 4378 3864 4380
rect 3888 4378 3944 4380
rect 3968 4378 4024 4380
rect 4048 4378 4104 4380
rect 3808 4326 3834 4378
rect 3834 4326 3864 4378
rect 3888 4326 3898 4378
rect 3898 4326 3944 4378
rect 3968 4326 4014 4378
rect 4014 4326 4024 4378
rect 4048 4326 4078 4378
rect 4078 4326 4104 4378
rect 3808 4324 3864 4326
rect 3888 4324 3944 4326
rect 3968 4324 4024 4326
rect 4048 4324 4104 4326
rect 3808 3290 3864 3292
rect 3888 3290 3944 3292
rect 3968 3290 4024 3292
rect 4048 3290 4104 3292
rect 3808 3238 3834 3290
rect 3834 3238 3864 3290
rect 3888 3238 3898 3290
rect 3898 3238 3944 3290
rect 3968 3238 4014 3290
rect 4014 3238 4024 3290
rect 4048 3238 4078 3290
rect 4078 3238 4104 3290
rect 3808 3236 3864 3238
rect 3888 3236 3944 3238
rect 3968 3236 4024 3238
rect 4048 3236 4104 3238
rect 3808 2202 3864 2204
rect 3888 2202 3944 2204
rect 3968 2202 4024 2204
rect 4048 2202 4104 2204
rect 3808 2150 3834 2202
rect 3834 2150 3864 2202
rect 3888 2150 3898 2202
rect 3898 2150 3944 2202
rect 3968 2150 4014 2202
rect 4014 2150 4024 2202
rect 4048 2150 4078 2202
rect 4078 2150 4104 2202
rect 3808 2148 3864 2150
rect 3888 2148 3944 2150
rect 3968 2148 4024 2150
rect 4048 2148 4104 2150
rect 4758 7098 4814 7100
rect 4838 7098 4894 7100
rect 4918 7098 4974 7100
rect 4998 7098 5054 7100
rect 4758 7046 4784 7098
rect 4784 7046 4814 7098
rect 4838 7046 4848 7098
rect 4848 7046 4894 7098
rect 4918 7046 4964 7098
rect 4964 7046 4974 7098
rect 4998 7046 5028 7098
rect 5028 7046 5054 7098
rect 4758 7044 4814 7046
rect 4838 7044 4894 7046
rect 4918 7044 4974 7046
rect 4998 7044 5054 7046
rect 4758 6010 4814 6012
rect 4838 6010 4894 6012
rect 4918 6010 4974 6012
rect 4998 6010 5054 6012
rect 4758 5958 4784 6010
rect 4784 5958 4814 6010
rect 4838 5958 4848 6010
rect 4848 5958 4894 6010
rect 4918 5958 4964 6010
rect 4964 5958 4974 6010
rect 4998 5958 5028 6010
rect 5028 5958 5054 6010
rect 4758 5956 4814 5958
rect 4838 5956 4894 5958
rect 4918 5956 4974 5958
rect 4998 5956 5054 5958
rect 5709 7642 5765 7644
rect 5789 7642 5845 7644
rect 5869 7642 5925 7644
rect 5949 7642 6005 7644
rect 5709 7590 5735 7642
rect 5735 7590 5765 7642
rect 5789 7590 5799 7642
rect 5799 7590 5845 7642
rect 5869 7590 5915 7642
rect 5915 7590 5925 7642
rect 5949 7590 5979 7642
rect 5979 7590 6005 7642
rect 5709 7588 5765 7590
rect 5789 7588 5845 7590
rect 5869 7588 5925 7590
rect 5949 7588 6005 7590
rect 4802 5772 4858 5808
rect 4802 5752 4804 5772
rect 4804 5752 4856 5772
rect 4856 5752 4858 5772
rect 4758 4922 4814 4924
rect 4838 4922 4894 4924
rect 4918 4922 4974 4924
rect 4998 4922 5054 4924
rect 4758 4870 4784 4922
rect 4784 4870 4814 4922
rect 4838 4870 4848 4922
rect 4848 4870 4894 4922
rect 4918 4870 4964 4922
rect 4964 4870 4974 4922
rect 4998 4870 5028 4922
rect 5028 4870 5054 4922
rect 4758 4868 4814 4870
rect 4838 4868 4894 4870
rect 4918 4868 4974 4870
rect 4998 4868 5054 4870
rect 4758 3834 4814 3836
rect 4838 3834 4894 3836
rect 4918 3834 4974 3836
rect 4998 3834 5054 3836
rect 4758 3782 4784 3834
rect 4784 3782 4814 3834
rect 4838 3782 4848 3834
rect 4848 3782 4894 3834
rect 4918 3782 4964 3834
rect 4964 3782 4974 3834
rect 4998 3782 5028 3834
rect 5028 3782 5054 3834
rect 4758 3780 4814 3782
rect 4838 3780 4894 3782
rect 4918 3780 4974 3782
rect 4998 3780 5054 3782
rect 5446 6160 5502 6216
rect 4434 2760 4490 2816
rect 4894 2916 4950 2952
rect 4894 2896 4896 2916
rect 4896 2896 4948 2916
rect 4948 2896 4950 2916
rect 4758 2746 4814 2748
rect 4838 2746 4894 2748
rect 4918 2746 4974 2748
rect 4998 2746 5054 2748
rect 4758 2694 4784 2746
rect 4784 2694 4814 2746
rect 4838 2694 4848 2746
rect 4848 2694 4894 2746
rect 4918 2694 4964 2746
rect 4964 2694 4974 2746
rect 4998 2694 5028 2746
rect 5028 2694 5054 2746
rect 4758 2692 4814 2694
rect 4838 2692 4894 2694
rect 4918 2692 4974 2694
rect 4998 2692 5054 2694
rect 5709 6554 5765 6556
rect 5789 6554 5845 6556
rect 5869 6554 5925 6556
rect 5949 6554 6005 6556
rect 5709 6502 5735 6554
rect 5735 6502 5765 6554
rect 5789 6502 5799 6554
rect 5799 6502 5845 6554
rect 5869 6502 5915 6554
rect 5915 6502 5925 6554
rect 5949 6502 5979 6554
rect 5979 6502 6005 6554
rect 5709 6500 5765 6502
rect 5789 6500 5845 6502
rect 5869 6500 5925 6502
rect 5949 6500 6005 6502
rect 5709 5466 5765 5468
rect 5789 5466 5845 5468
rect 5869 5466 5925 5468
rect 5949 5466 6005 5468
rect 5709 5414 5735 5466
rect 5735 5414 5765 5466
rect 5789 5414 5799 5466
rect 5799 5414 5845 5466
rect 5869 5414 5915 5466
rect 5915 5414 5925 5466
rect 5949 5414 5979 5466
rect 5979 5414 6005 5466
rect 5709 5412 5765 5414
rect 5789 5412 5845 5414
rect 5869 5412 5925 5414
rect 5949 5412 6005 5414
rect 5709 4378 5765 4380
rect 5789 4378 5845 4380
rect 5869 4378 5925 4380
rect 5949 4378 6005 4380
rect 5709 4326 5735 4378
rect 5735 4326 5765 4378
rect 5789 4326 5799 4378
rect 5799 4326 5845 4378
rect 5869 4326 5915 4378
rect 5915 4326 5925 4378
rect 5949 4326 5979 4378
rect 5979 4326 6005 4378
rect 5709 4324 5765 4326
rect 5789 4324 5845 4326
rect 5869 4324 5925 4326
rect 5949 4324 6005 4326
rect 6090 3440 6146 3496
rect 5709 3290 5765 3292
rect 5789 3290 5845 3292
rect 5869 3290 5925 3292
rect 5949 3290 6005 3292
rect 5709 3238 5735 3290
rect 5735 3238 5765 3290
rect 5789 3238 5799 3290
rect 5799 3238 5845 3290
rect 5869 3238 5915 3290
rect 5915 3238 5925 3290
rect 5949 3238 5979 3290
rect 5979 3238 6005 3290
rect 5709 3236 5765 3238
rect 5789 3236 5845 3238
rect 5869 3236 5925 3238
rect 5949 3236 6005 3238
rect 5709 2202 5765 2204
rect 5789 2202 5845 2204
rect 5869 2202 5925 2204
rect 5949 2202 6005 2204
rect 5709 2150 5735 2202
rect 5735 2150 5765 2202
rect 5789 2150 5799 2202
rect 5799 2150 5845 2202
rect 5869 2150 5915 2202
rect 5915 2150 5925 2202
rect 5949 2150 5979 2202
rect 5979 2150 6005 2202
rect 5709 2148 5765 2150
rect 5789 2148 5845 2150
rect 5869 2148 5925 2150
rect 5949 2148 6005 2150
rect 3698 720 3754 776
<< metal3 >>
rect 0 8938 800 8968
rect 2773 8938 2839 8941
rect 0 8936 2839 8938
rect 0 8880 2778 8936
rect 2834 8880 2839 8936
rect 0 8878 2839 8880
rect 0 8848 800 8878
rect 2773 8875 2839 8878
rect 1894 7648 2214 7649
rect 1894 7584 1902 7648
rect 1966 7584 1982 7648
rect 2046 7584 2062 7648
rect 2126 7584 2142 7648
rect 2206 7584 2214 7648
rect 1894 7583 2214 7584
rect 3796 7648 4116 7649
rect 3796 7584 3804 7648
rect 3868 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4116 7648
rect 3796 7583 4116 7584
rect 5697 7648 6017 7649
rect 5697 7584 5705 7648
rect 5769 7584 5785 7648
rect 5849 7584 5865 7648
rect 5929 7584 5945 7648
rect 6009 7584 6017 7648
rect 5697 7583 6017 7584
rect 2845 7104 3165 7105
rect 2845 7040 2853 7104
rect 2917 7040 2933 7104
rect 2997 7040 3013 7104
rect 3077 7040 3093 7104
rect 3157 7040 3165 7104
rect 2845 7039 3165 7040
rect 4746 7104 5066 7105
rect 4746 7040 4754 7104
rect 4818 7040 4834 7104
rect 4898 7040 4914 7104
rect 4978 7040 4994 7104
rect 5058 7040 5066 7104
rect 4746 7039 5066 7040
rect 1894 6560 2214 6561
rect 1894 6496 1902 6560
rect 1966 6496 1982 6560
rect 2046 6496 2062 6560
rect 2126 6496 2142 6560
rect 2206 6496 2214 6560
rect 1894 6495 2214 6496
rect 3796 6560 4116 6561
rect 3796 6496 3804 6560
rect 3868 6496 3884 6560
rect 3948 6496 3964 6560
rect 4028 6496 4044 6560
rect 4108 6496 4116 6560
rect 3796 6495 4116 6496
rect 5697 6560 6017 6561
rect 5697 6496 5705 6560
rect 5769 6496 5785 6560
rect 5849 6496 5865 6560
rect 5929 6496 5945 6560
rect 6009 6496 6017 6560
rect 5697 6495 6017 6496
rect 0 6218 800 6248
rect 1761 6218 1827 6221
rect 0 6216 1827 6218
rect 0 6160 1766 6216
rect 1822 6160 1827 6216
rect 0 6158 1827 6160
rect 0 6128 800 6158
rect 1761 6155 1827 6158
rect 5441 6218 5507 6221
rect 7199 6218 7999 6248
rect 5441 6216 7999 6218
rect 5441 6160 5446 6216
rect 5502 6160 7999 6216
rect 5441 6158 7999 6160
rect 5441 6155 5507 6158
rect 7199 6128 7999 6158
rect 2845 6016 3165 6017
rect 2845 5952 2853 6016
rect 2917 5952 2933 6016
rect 2997 5952 3013 6016
rect 3077 5952 3093 6016
rect 3157 5952 3165 6016
rect 2845 5951 3165 5952
rect 4746 6016 5066 6017
rect 4746 5952 4754 6016
rect 4818 5952 4834 6016
rect 4898 5952 4914 6016
rect 4978 5952 4994 6016
rect 5058 5952 5066 6016
rect 4746 5951 5066 5952
rect 3233 5810 3299 5813
rect 4245 5810 4311 5813
rect 4797 5810 4863 5813
rect 3233 5808 4863 5810
rect 3233 5752 3238 5808
rect 3294 5752 4250 5808
rect 4306 5752 4802 5808
rect 4858 5752 4863 5808
rect 3233 5750 4863 5752
rect 3233 5747 3299 5750
rect 4245 5747 4311 5750
rect 4797 5747 4863 5750
rect 1894 5472 2214 5473
rect 1894 5408 1902 5472
rect 1966 5408 1982 5472
rect 2046 5408 2062 5472
rect 2126 5408 2142 5472
rect 2206 5408 2214 5472
rect 1894 5407 2214 5408
rect 3796 5472 4116 5473
rect 3796 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4116 5472
rect 3796 5407 4116 5408
rect 5697 5472 6017 5473
rect 5697 5408 5705 5472
rect 5769 5408 5785 5472
rect 5849 5408 5865 5472
rect 5929 5408 5945 5472
rect 6009 5408 6017 5472
rect 5697 5407 6017 5408
rect 2845 4928 3165 4929
rect 2845 4864 2853 4928
rect 2917 4864 2933 4928
rect 2997 4864 3013 4928
rect 3077 4864 3093 4928
rect 3157 4864 3165 4928
rect 2845 4863 3165 4864
rect 4746 4928 5066 4929
rect 4746 4864 4754 4928
rect 4818 4864 4834 4928
rect 4898 4864 4914 4928
rect 4978 4864 4994 4928
rect 5058 4864 5066 4928
rect 4746 4863 5066 4864
rect 1894 4384 2214 4385
rect 1894 4320 1902 4384
rect 1966 4320 1982 4384
rect 2046 4320 2062 4384
rect 2126 4320 2142 4384
rect 2206 4320 2214 4384
rect 1894 4319 2214 4320
rect 3796 4384 4116 4385
rect 3796 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4116 4384
rect 3796 4319 4116 4320
rect 5697 4384 6017 4385
rect 5697 4320 5705 4384
rect 5769 4320 5785 4384
rect 5849 4320 5865 4384
rect 5929 4320 5945 4384
rect 6009 4320 6017 4384
rect 5697 4319 6017 4320
rect 2845 3840 3165 3841
rect 2845 3776 2853 3840
rect 2917 3776 2933 3840
rect 2997 3776 3013 3840
rect 3077 3776 3093 3840
rect 3157 3776 3165 3840
rect 2845 3775 3165 3776
rect 4746 3840 5066 3841
rect 4746 3776 4754 3840
rect 4818 3776 4834 3840
rect 4898 3776 4914 3840
rect 4978 3776 4994 3840
rect 5058 3776 5066 3840
rect 4746 3775 5066 3776
rect 0 3498 800 3528
rect 1761 3498 1827 3501
rect 0 3496 1827 3498
rect 0 3440 1766 3496
rect 1822 3440 1827 3496
rect 0 3438 1827 3440
rect 0 3408 800 3438
rect 1761 3435 1827 3438
rect 6085 3498 6151 3501
rect 7199 3498 7999 3528
rect 6085 3496 7999 3498
rect 6085 3440 6090 3496
rect 6146 3440 7999 3496
rect 6085 3438 7999 3440
rect 6085 3435 6151 3438
rect 7199 3408 7999 3438
rect 1894 3296 2214 3297
rect 1894 3232 1902 3296
rect 1966 3232 1982 3296
rect 2046 3232 2062 3296
rect 2126 3232 2142 3296
rect 2206 3232 2214 3296
rect 1894 3231 2214 3232
rect 3796 3296 4116 3297
rect 3796 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4116 3296
rect 3796 3231 4116 3232
rect 5697 3296 6017 3297
rect 5697 3232 5705 3296
rect 5769 3232 5785 3296
rect 5849 3232 5865 3296
rect 5929 3232 5945 3296
rect 6009 3232 6017 3296
rect 5697 3231 6017 3232
rect 4889 2954 4955 2957
rect 4478 2952 4955 2954
rect 4478 2896 4894 2952
rect 4950 2896 4955 2952
rect 4478 2894 4955 2896
rect 4478 2821 4538 2894
rect 4889 2891 4955 2894
rect 4429 2816 4538 2821
rect 4429 2760 4434 2816
rect 4490 2760 4538 2816
rect 4429 2758 4538 2760
rect 4429 2755 4495 2758
rect 2845 2752 3165 2753
rect 2845 2688 2853 2752
rect 2917 2688 2933 2752
rect 2997 2688 3013 2752
rect 3077 2688 3093 2752
rect 3157 2688 3165 2752
rect 2845 2687 3165 2688
rect 4746 2752 5066 2753
rect 4746 2688 4754 2752
rect 4818 2688 4834 2752
rect 4898 2688 4914 2752
rect 4978 2688 4994 2752
rect 5058 2688 5066 2752
rect 4746 2687 5066 2688
rect 1894 2208 2214 2209
rect 1894 2144 1902 2208
rect 1966 2144 1982 2208
rect 2046 2144 2062 2208
rect 2126 2144 2142 2208
rect 2206 2144 2214 2208
rect 1894 2143 2214 2144
rect 3796 2208 4116 2209
rect 3796 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4116 2208
rect 3796 2143 4116 2144
rect 5697 2208 6017 2209
rect 5697 2144 5705 2208
rect 5769 2144 5785 2208
rect 5849 2144 5865 2208
rect 5929 2144 5945 2208
rect 6009 2144 6017 2208
rect 5697 2143 6017 2144
rect 3693 778 3759 781
rect 7199 778 7999 808
rect 3693 776 7999 778
rect 3693 720 3698 776
rect 3754 720 7999 776
rect 3693 718 7999 720
rect 3693 715 3759 718
rect 7199 688 7999 718
<< via3 >>
rect 1902 7644 1966 7648
rect 1902 7588 1906 7644
rect 1906 7588 1962 7644
rect 1962 7588 1966 7644
rect 1902 7584 1966 7588
rect 1982 7644 2046 7648
rect 1982 7588 1986 7644
rect 1986 7588 2042 7644
rect 2042 7588 2046 7644
rect 1982 7584 2046 7588
rect 2062 7644 2126 7648
rect 2062 7588 2066 7644
rect 2066 7588 2122 7644
rect 2122 7588 2126 7644
rect 2062 7584 2126 7588
rect 2142 7644 2206 7648
rect 2142 7588 2146 7644
rect 2146 7588 2202 7644
rect 2202 7588 2206 7644
rect 2142 7584 2206 7588
rect 3804 7644 3868 7648
rect 3804 7588 3808 7644
rect 3808 7588 3864 7644
rect 3864 7588 3868 7644
rect 3804 7584 3868 7588
rect 3884 7644 3948 7648
rect 3884 7588 3888 7644
rect 3888 7588 3944 7644
rect 3944 7588 3948 7644
rect 3884 7584 3948 7588
rect 3964 7644 4028 7648
rect 3964 7588 3968 7644
rect 3968 7588 4024 7644
rect 4024 7588 4028 7644
rect 3964 7584 4028 7588
rect 4044 7644 4108 7648
rect 4044 7588 4048 7644
rect 4048 7588 4104 7644
rect 4104 7588 4108 7644
rect 4044 7584 4108 7588
rect 5705 7644 5769 7648
rect 5705 7588 5709 7644
rect 5709 7588 5765 7644
rect 5765 7588 5769 7644
rect 5705 7584 5769 7588
rect 5785 7644 5849 7648
rect 5785 7588 5789 7644
rect 5789 7588 5845 7644
rect 5845 7588 5849 7644
rect 5785 7584 5849 7588
rect 5865 7644 5929 7648
rect 5865 7588 5869 7644
rect 5869 7588 5925 7644
rect 5925 7588 5929 7644
rect 5865 7584 5929 7588
rect 5945 7644 6009 7648
rect 5945 7588 5949 7644
rect 5949 7588 6005 7644
rect 6005 7588 6009 7644
rect 5945 7584 6009 7588
rect 2853 7100 2917 7104
rect 2853 7044 2857 7100
rect 2857 7044 2913 7100
rect 2913 7044 2917 7100
rect 2853 7040 2917 7044
rect 2933 7100 2997 7104
rect 2933 7044 2937 7100
rect 2937 7044 2993 7100
rect 2993 7044 2997 7100
rect 2933 7040 2997 7044
rect 3013 7100 3077 7104
rect 3013 7044 3017 7100
rect 3017 7044 3073 7100
rect 3073 7044 3077 7100
rect 3013 7040 3077 7044
rect 3093 7100 3157 7104
rect 3093 7044 3097 7100
rect 3097 7044 3153 7100
rect 3153 7044 3157 7100
rect 3093 7040 3157 7044
rect 4754 7100 4818 7104
rect 4754 7044 4758 7100
rect 4758 7044 4814 7100
rect 4814 7044 4818 7100
rect 4754 7040 4818 7044
rect 4834 7100 4898 7104
rect 4834 7044 4838 7100
rect 4838 7044 4894 7100
rect 4894 7044 4898 7100
rect 4834 7040 4898 7044
rect 4914 7100 4978 7104
rect 4914 7044 4918 7100
rect 4918 7044 4974 7100
rect 4974 7044 4978 7100
rect 4914 7040 4978 7044
rect 4994 7100 5058 7104
rect 4994 7044 4998 7100
rect 4998 7044 5054 7100
rect 5054 7044 5058 7100
rect 4994 7040 5058 7044
rect 1902 6556 1966 6560
rect 1902 6500 1906 6556
rect 1906 6500 1962 6556
rect 1962 6500 1966 6556
rect 1902 6496 1966 6500
rect 1982 6556 2046 6560
rect 1982 6500 1986 6556
rect 1986 6500 2042 6556
rect 2042 6500 2046 6556
rect 1982 6496 2046 6500
rect 2062 6556 2126 6560
rect 2062 6500 2066 6556
rect 2066 6500 2122 6556
rect 2122 6500 2126 6556
rect 2062 6496 2126 6500
rect 2142 6556 2206 6560
rect 2142 6500 2146 6556
rect 2146 6500 2202 6556
rect 2202 6500 2206 6556
rect 2142 6496 2206 6500
rect 3804 6556 3868 6560
rect 3804 6500 3808 6556
rect 3808 6500 3864 6556
rect 3864 6500 3868 6556
rect 3804 6496 3868 6500
rect 3884 6556 3948 6560
rect 3884 6500 3888 6556
rect 3888 6500 3944 6556
rect 3944 6500 3948 6556
rect 3884 6496 3948 6500
rect 3964 6556 4028 6560
rect 3964 6500 3968 6556
rect 3968 6500 4024 6556
rect 4024 6500 4028 6556
rect 3964 6496 4028 6500
rect 4044 6556 4108 6560
rect 4044 6500 4048 6556
rect 4048 6500 4104 6556
rect 4104 6500 4108 6556
rect 4044 6496 4108 6500
rect 5705 6556 5769 6560
rect 5705 6500 5709 6556
rect 5709 6500 5765 6556
rect 5765 6500 5769 6556
rect 5705 6496 5769 6500
rect 5785 6556 5849 6560
rect 5785 6500 5789 6556
rect 5789 6500 5845 6556
rect 5845 6500 5849 6556
rect 5785 6496 5849 6500
rect 5865 6556 5929 6560
rect 5865 6500 5869 6556
rect 5869 6500 5925 6556
rect 5925 6500 5929 6556
rect 5865 6496 5929 6500
rect 5945 6556 6009 6560
rect 5945 6500 5949 6556
rect 5949 6500 6005 6556
rect 6005 6500 6009 6556
rect 5945 6496 6009 6500
rect 2853 6012 2917 6016
rect 2853 5956 2857 6012
rect 2857 5956 2913 6012
rect 2913 5956 2917 6012
rect 2853 5952 2917 5956
rect 2933 6012 2997 6016
rect 2933 5956 2937 6012
rect 2937 5956 2993 6012
rect 2993 5956 2997 6012
rect 2933 5952 2997 5956
rect 3013 6012 3077 6016
rect 3013 5956 3017 6012
rect 3017 5956 3073 6012
rect 3073 5956 3077 6012
rect 3013 5952 3077 5956
rect 3093 6012 3157 6016
rect 3093 5956 3097 6012
rect 3097 5956 3153 6012
rect 3153 5956 3157 6012
rect 3093 5952 3157 5956
rect 4754 6012 4818 6016
rect 4754 5956 4758 6012
rect 4758 5956 4814 6012
rect 4814 5956 4818 6012
rect 4754 5952 4818 5956
rect 4834 6012 4898 6016
rect 4834 5956 4838 6012
rect 4838 5956 4894 6012
rect 4894 5956 4898 6012
rect 4834 5952 4898 5956
rect 4914 6012 4978 6016
rect 4914 5956 4918 6012
rect 4918 5956 4974 6012
rect 4974 5956 4978 6012
rect 4914 5952 4978 5956
rect 4994 6012 5058 6016
rect 4994 5956 4998 6012
rect 4998 5956 5054 6012
rect 5054 5956 5058 6012
rect 4994 5952 5058 5956
rect 1902 5468 1966 5472
rect 1902 5412 1906 5468
rect 1906 5412 1962 5468
rect 1962 5412 1966 5468
rect 1902 5408 1966 5412
rect 1982 5468 2046 5472
rect 1982 5412 1986 5468
rect 1986 5412 2042 5468
rect 2042 5412 2046 5468
rect 1982 5408 2046 5412
rect 2062 5468 2126 5472
rect 2062 5412 2066 5468
rect 2066 5412 2122 5468
rect 2122 5412 2126 5468
rect 2062 5408 2126 5412
rect 2142 5468 2206 5472
rect 2142 5412 2146 5468
rect 2146 5412 2202 5468
rect 2202 5412 2206 5468
rect 2142 5408 2206 5412
rect 3804 5468 3868 5472
rect 3804 5412 3808 5468
rect 3808 5412 3864 5468
rect 3864 5412 3868 5468
rect 3804 5408 3868 5412
rect 3884 5468 3948 5472
rect 3884 5412 3888 5468
rect 3888 5412 3944 5468
rect 3944 5412 3948 5468
rect 3884 5408 3948 5412
rect 3964 5468 4028 5472
rect 3964 5412 3968 5468
rect 3968 5412 4024 5468
rect 4024 5412 4028 5468
rect 3964 5408 4028 5412
rect 4044 5468 4108 5472
rect 4044 5412 4048 5468
rect 4048 5412 4104 5468
rect 4104 5412 4108 5468
rect 4044 5408 4108 5412
rect 5705 5468 5769 5472
rect 5705 5412 5709 5468
rect 5709 5412 5765 5468
rect 5765 5412 5769 5468
rect 5705 5408 5769 5412
rect 5785 5468 5849 5472
rect 5785 5412 5789 5468
rect 5789 5412 5845 5468
rect 5845 5412 5849 5468
rect 5785 5408 5849 5412
rect 5865 5468 5929 5472
rect 5865 5412 5869 5468
rect 5869 5412 5925 5468
rect 5925 5412 5929 5468
rect 5865 5408 5929 5412
rect 5945 5468 6009 5472
rect 5945 5412 5949 5468
rect 5949 5412 6005 5468
rect 6005 5412 6009 5468
rect 5945 5408 6009 5412
rect 2853 4924 2917 4928
rect 2853 4868 2857 4924
rect 2857 4868 2913 4924
rect 2913 4868 2917 4924
rect 2853 4864 2917 4868
rect 2933 4924 2997 4928
rect 2933 4868 2937 4924
rect 2937 4868 2993 4924
rect 2993 4868 2997 4924
rect 2933 4864 2997 4868
rect 3013 4924 3077 4928
rect 3013 4868 3017 4924
rect 3017 4868 3073 4924
rect 3073 4868 3077 4924
rect 3013 4864 3077 4868
rect 3093 4924 3157 4928
rect 3093 4868 3097 4924
rect 3097 4868 3153 4924
rect 3153 4868 3157 4924
rect 3093 4864 3157 4868
rect 4754 4924 4818 4928
rect 4754 4868 4758 4924
rect 4758 4868 4814 4924
rect 4814 4868 4818 4924
rect 4754 4864 4818 4868
rect 4834 4924 4898 4928
rect 4834 4868 4838 4924
rect 4838 4868 4894 4924
rect 4894 4868 4898 4924
rect 4834 4864 4898 4868
rect 4914 4924 4978 4928
rect 4914 4868 4918 4924
rect 4918 4868 4974 4924
rect 4974 4868 4978 4924
rect 4914 4864 4978 4868
rect 4994 4924 5058 4928
rect 4994 4868 4998 4924
rect 4998 4868 5054 4924
rect 5054 4868 5058 4924
rect 4994 4864 5058 4868
rect 1902 4380 1966 4384
rect 1902 4324 1906 4380
rect 1906 4324 1962 4380
rect 1962 4324 1966 4380
rect 1902 4320 1966 4324
rect 1982 4380 2046 4384
rect 1982 4324 1986 4380
rect 1986 4324 2042 4380
rect 2042 4324 2046 4380
rect 1982 4320 2046 4324
rect 2062 4380 2126 4384
rect 2062 4324 2066 4380
rect 2066 4324 2122 4380
rect 2122 4324 2126 4380
rect 2062 4320 2126 4324
rect 2142 4380 2206 4384
rect 2142 4324 2146 4380
rect 2146 4324 2202 4380
rect 2202 4324 2206 4380
rect 2142 4320 2206 4324
rect 3804 4380 3868 4384
rect 3804 4324 3808 4380
rect 3808 4324 3864 4380
rect 3864 4324 3868 4380
rect 3804 4320 3868 4324
rect 3884 4380 3948 4384
rect 3884 4324 3888 4380
rect 3888 4324 3944 4380
rect 3944 4324 3948 4380
rect 3884 4320 3948 4324
rect 3964 4380 4028 4384
rect 3964 4324 3968 4380
rect 3968 4324 4024 4380
rect 4024 4324 4028 4380
rect 3964 4320 4028 4324
rect 4044 4380 4108 4384
rect 4044 4324 4048 4380
rect 4048 4324 4104 4380
rect 4104 4324 4108 4380
rect 4044 4320 4108 4324
rect 5705 4380 5769 4384
rect 5705 4324 5709 4380
rect 5709 4324 5765 4380
rect 5765 4324 5769 4380
rect 5705 4320 5769 4324
rect 5785 4380 5849 4384
rect 5785 4324 5789 4380
rect 5789 4324 5845 4380
rect 5845 4324 5849 4380
rect 5785 4320 5849 4324
rect 5865 4380 5929 4384
rect 5865 4324 5869 4380
rect 5869 4324 5925 4380
rect 5925 4324 5929 4380
rect 5865 4320 5929 4324
rect 5945 4380 6009 4384
rect 5945 4324 5949 4380
rect 5949 4324 6005 4380
rect 6005 4324 6009 4380
rect 5945 4320 6009 4324
rect 2853 3836 2917 3840
rect 2853 3780 2857 3836
rect 2857 3780 2913 3836
rect 2913 3780 2917 3836
rect 2853 3776 2917 3780
rect 2933 3836 2997 3840
rect 2933 3780 2937 3836
rect 2937 3780 2993 3836
rect 2993 3780 2997 3836
rect 2933 3776 2997 3780
rect 3013 3836 3077 3840
rect 3013 3780 3017 3836
rect 3017 3780 3073 3836
rect 3073 3780 3077 3836
rect 3013 3776 3077 3780
rect 3093 3836 3157 3840
rect 3093 3780 3097 3836
rect 3097 3780 3153 3836
rect 3153 3780 3157 3836
rect 3093 3776 3157 3780
rect 4754 3836 4818 3840
rect 4754 3780 4758 3836
rect 4758 3780 4814 3836
rect 4814 3780 4818 3836
rect 4754 3776 4818 3780
rect 4834 3836 4898 3840
rect 4834 3780 4838 3836
rect 4838 3780 4894 3836
rect 4894 3780 4898 3836
rect 4834 3776 4898 3780
rect 4914 3836 4978 3840
rect 4914 3780 4918 3836
rect 4918 3780 4974 3836
rect 4974 3780 4978 3836
rect 4914 3776 4978 3780
rect 4994 3836 5058 3840
rect 4994 3780 4998 3836
rect 4998 3780 5054 3836
rect 5054 3780 5058 3836
rect 4994 3776 5058 3780
rect 1902 3292 1966 3296
rect 1902 3236 1906 3292
rect 1906 3236 1962 3292
rect 1962 3236 1966 3292
rect 1902 3232 1966 3236
rect 1982 3292 2046 3296
rect 1982 3236 1986 3292
rect 1986 3236 2042 3292
rect 2042 3236 2046 3292
rect 1982 3232 2046 3236
rect 2062 3292 2126 3296
rect 2062 3236 2066 3292
rect 2066 3236 2122 3292
rect 2122 3236 2126 3292
rect 2062 3232 2126 3236
rect 2142 3292 2206 3296
rect 2142 3236 2146 3292
rect 2146 3236 2202 3292
rect 2202 3236 2206 3292
rect 2142 3232 2206 3236
rect 3804 3292 3868 3296
rect 3804 3236 3808 3292
rect 3808 3236 3864 3292
rect 3864 3236 3868 3292
rect 3804 3232 3868 3236
rect 3884 3292 3948 3296
rect 3884 3236 3888 3292
rect 3888 3236 3944 3292
rect 3944 3236 3948 3292
rect 3884 3232 3948 3236
rect 3964 3292 4028 3296
rect 3964 3236 3968 3292
rect 3968 3236 4024 3292
rect 4024 3236 4028 3292
rect 3964 3232 4028 3236
rect 4044 3292 4108 3296
rect 4044 3236 4048 3292
rect 4048 3236 4104 3292
rect 4104 3236 4108 3292
rect 4044 3232 4108 3236
rect 5705 3292 5769 3296
rect 5705 3236 5709 3292
rect 5709 3236 5765 3292
rect 5765 3236 5769 3292
rect 5705 3232 5769 3236
rect 5785 3292 5849 3296
rect 5785 3236 5789 3292
rect 5789 3236 5845 3292
rect 5845 3236 5849 3292
rect 5785 3232 5849 3236
rect 5865 3292 5929 3296
rect 5865 3236 5869 3292
rect 5869 3236 5925 3292
rect 5925 3236 5929 3292
rect 5865 3232 5929 3236
rect 5945 3292 6009 3296
rect 5945 3236 5949 3292
rect 5949 3236 6005 3292
rect 6005 3236 6009 3292
rect 5945 3232 6009 3236
rect 2853 2748 2917 2752
rect 2853 2692 2857 2748
rect 2857 2692 2913 2748
rect 2913 2692 2917 2748
rect 2853 2688 2917 2692
rect 2933 2748 2997 2752
rect 2933 2692 2937 2748
rect 2937 2692 2993 2748
rect 2993 2692 2997 2748
rect 2933 2688 2997 2692
rect 3013 2748 3077 2752
rect 3013 2692 3017 2748
rect 3017 2692 3073 2748
rect 3073 2692 3077 2748
rect 3013 2688 3077 2692
rect 3093 2748 3157 2752
rect 3093 2692 3097 2748
rect 3097 2692 3153 2748
rect 3153 2692 3157 2748
rect 3093 2688 3157 2692
rect 4754 2748 4818 2752
rect 4754 2692 4758 2748
rect 4758 2692 4814 2748
rect 4814 2692 4818 2748
rect 4754 2688 4818 2692
rect 4834 2748 4898 2752
rect 4834 2692 4838 2748
rect 4838 2692 4894 2748
rect 4894 2692 4898 2748
rect 4834 2688 4898 2692
rect 4914 2748 4978 2752
rect 4914 2692 4918 2748
rect 4918 2692 4974 2748
rect 4974 2692 4978 2748
rect 4914 2688 4978 2692
rect 4994 2748 5058 2752
rect 4994 2692 4998 2748
rect 4998 2692 5054 2748
rect 5054 2692 5058 2748
rect 4994 2688 5058 2692
rect 1902 2204 1966 2208
rect 1902 2148 1906 2204
rect 1906 2148 1962 2204
rect 1962 2148 1966 2204
rect 1902 2144 1966 2148
rect 1982 2204 2046 2208
rect 1982 2148 1986 2204
rect 1986 2148 2042 2204
rect 2042 2148 2046 2204
rect 1982 2144 2046 2148
rect 2062 2204 2126 2208
rect 2062 2148 2066 2204
rect 2066 2148 2122 2204
rect 2122 2148 2126 2204
rect 2062 2144 2126 2148
rect 2142 2204 2206 2208
rect 2142 2148 2146 2204
rect 2146 2148 2202 2204
rect 2202 2148 2206 2204
rect 2142 2144 2206 2148
rect 3804 2204 3868 2208
rect 3804 2148 3808 2204
rect 3808 2148 3864 2204
rect 3864 2148 3868 2204
rect 3804 2144 3868 2148
rect 3884 2204 3948 2208
rect 3884 2148 3888 2204
rect 3888 2148 3944 2204
rect 3944 2148 3948 2204
rect 3884 2144 3948 2148
rect 3964 2204 4028 2208
rect 3964 2148 3968 2204
rect 3968 2148 4024 2204
rect 4024 2148 4028 2204
rect 3964 2144 4028 2148
rect 4044 2204 4108 2208
rect 4044 2148 4048 2204
rect 4048 2148 4104 2204
rect 4104 2148 4108 2204
rect 4044 2144 4108 2148
rect 5705 2204 5769 2208
rect 5705 2148 5709 2204
rect 5709 2148 5765 2204
rect 5765 2148 5769 2204
rect 5705 2144 5769 2148
rect 5785 2204 5849 2208
rect 5785 2148 5789 2204
rect 5789 2148 5845 2204
rect 5845 2148 5849 2204
rect 5785 2144 5849 2148
rect 5865 2204 5929 2208
rect 5865 2148 5869 2204
rect 5869 2148 5925 2204
rect 5925 2148 5929 2204
rect 5865 2144 5929 2148
rect 5945 2204 6009 2208
rect 5945 2148 5949 2204
rect 5949 2148 6005 2204
rect 6005 2148 6009 2204
rect 5945 2144 6009 2148
<< metal4 >>
rect 1894 7648 2215 7664
rect 1894 7584 1902 7648
rect 1966 7584 1982 7648
rect 2046 7584 2062 7648
rect 2126 7584 2142 7648
rect 2206 7584 2215 7648
rect 1894 6779 2215 7584
rect 1894 6560 1936 6779
rect 2172 6560 2215 6779
rect 1894 6496 1902 6560
rect 1966 6496 1982 6543
rect 2046 6496 2062 6543
rect 2126 6496 2142 6543
rect 2206 6496 2215 6560
rect 1894 5472 2215 6496
rect 1894 5408 1902 5472
rect 1966 5408 1982 5472
rect 2046 5408 2062 5472
rect 2126 5408 2142 5472
rect 2206 5408 2215 5472
rect 1894 4966 2215 5408
rect 1894 4730 1936 4966
rect 2172 4730 2215 4966
rect 1894 4384 2215 4730
rect 1894 4320 1902 4384
rect 1966 4320 1982 4384
rect 2046 4320 2062 4384
rect 2126 4320 2142 4384
rect 2206 4320 2215 4384
rect 1894 3296 2215 4320
rect 1894 3232 1902 3296
rect 1966 3232 1982 3296
rect 2046 3232 2062 3296
rect 2126 3232 2142 3296
rect 2206 3232 2215 3296
rect 1894 3152 2215 3232
rect 1894 2916 1936 3152
rect 2172 2916 2215 3152
rect 1894 2208 2215 2916
rect 1894 2144 1902 2208
rect 1966 2144 1982 2208
rect 2046 2144 2062 2208
rect 2126 2144 2142 2208
rect 2206 2144 2215 2208
rect 1894 2128 2215 2144
rect 2845 7104 3165 7664
rect 2845 7040 2853 7104
rect 2917 7040 2933 7104
rect 2997 7040 3013 7104
rect 3077 7040 3093 7104
rect 3157 7040 3165 7104
rect 2845 6016 3165 7040
rect 2845 5952 2853 6016
rect 2917 5952 2933 6016
rect 2997 5952 3013 6016
rect 3077 5952 3093 6016
rect 3157 5952 3165 6016
rect 2845 5872 3165 5952
rect 2845 5636 2887 5872
rect 3123 5636 3165 5872
rect 2845 4928 3165 5636
rect 2845 4864 2853 4928
rect 2917 4864 2933 4928
rect 2997 4864 3013 4928
rect 3077 4864 3093 4928
rect 3157 4864 3165 4928
rect 2845 4059 3165 4864
rect 2845 3840 2887 4059
rect 3123 3840 3165 4059
rect 2845 3776 2853 3840
rect 2917 3776 2933 3823
rect 2997 3776 3013 3823
rect 3077 3776 3093 3823
rect 3157 3776 3165 3840
rect 2845 2752 3165 3776
rect 2845 2688 2853 2752
rect 2917 2688 2933 2752
rect 2997 2688 3013 2752
rect 3077 2688 3093 2752
rect 3157 2688 3165 2752
rect 2845 2128 3165 2688
rect 3796 7648 4116 7664
rect 3796 7584 3804 7648
rect 3868 7584 3884 7648
rect 3948 7584 3964 7648
rect 4028 7584 4044 7648
rect 4108 7584 4116 7648
rect 3796 6779 4116 7584
rect 3796 6560 3838 6779
rect 4074 6560 4116 6779
rect 3796 6496 3804 6560
rect 3868 6496 3884 6543
rect 3948 6496 3964 6543
rect 4028 6496 4044 6543
rect 4108 6496 4116 6560
rect 3796 5472 4116 6496
rect 3796 5408 3804 5472
rect 3868 5408 3884 5472
rect 3948 5408 3964 5472
rect 4028 5408 4044 5472
rect 4108 5408 4116 5472
rect 3796 4966 4116 5408
rect 3796 4730 3838 4966
rect 4074 4730 4116 4966
rect 3796 4384 4116 4730
rect 3796 4320 3804 4384
rect 3868 4320 3884 4384
rect 3948 4320 3964 4384
rect 4028 4320 4044 4384
rect 4108 4320 4116 4384
rect 3796 3296 4116 4320
rect 3796 3232 3804 3296
rect 3868 3232 3884 3296
rect 3948 3232 3964 3296
rect 4028 3232 4044 3296
rect 4108 3232 4116 3296
rect 3796 3152 4116 3232
rect 3796 2916 3838 3152
rect 4074 2916 4116 3152
rect 3796 2208 4116 2916
rect 3796 2144 3804 2208
rect 3868 2144 3884 2208
rect 3948 2144 3964 2208
rect 4028 2144 4044 2208
rect 4108 2144 4116 2208
rect 3796 2128 4116 2144
rect 4746 7104 5067 7664
rect 4746 7040 4754 7104
rect 4818 7040 4834 7104
rect 4898 7040 4914 7104
rect 4978 7040 4994 7104
rect 5058 7040 5067 7104
rect 4746 6016 5067 7040
rect 4746 5952 4754 6016
rect 4818 5952 4834 6016
rect 4898 5952 4914 6016
rect 4978 5952 4994 6016
rect 5058 5952 5067 6016
rect 4746 5872 5067 5952
rect 4746 5636 4788 5872
rect 5024 5636 5067 5872
rect 4746 4928 5067 5636
rect 4746 4864 4754 4928
rect 4818 4864 4834 4928
rect 4898 4864 4914 4928
rect 4978 4864 4994 4928
rect 5058 4864 5067 4928
rect 4746 4059 5067 4864
rect 4746 3840 4788 4059
rect 5024 3840 5067 4059
rect 4746 3776 4754 3840
rect 4818 3776 4834 3823
rect 4898 3776 4914 3823
rect 4978 3776 4994 3823
rect 5058 3776 5067 3840
rect 4746 2752 5067 3776
rect 4746 2688 4754 2752
rect 4818 2688 4834 2752
rect 4898 2688 4914 2752
rect 4978 2688 4994 2752
rect 5058 2688 5067 2752
rect 4746 2128 5067 2688
rect 5697 7648 6017 7664
rect 5697 7584 5705 7648
rect 5769 7584 5785 7648
rect 5849 7584 5865 7648
rect 5929 7584 5945 7648
rect 6009 7584 6017 7648
rect 5697 6779 6017 7584
rect 5697 6560 5739 6779
rect 5975 6560 6017 6779
rect 5697 6496 5705 6560
rect 5769 6496 5785 6543
rect 5849 6496 5865 6543
rect 5929 6496 5945 6543
rect 6009 6496 6017 6560
rect 5697 5472 6017 6496
rect 5697 5408 5705 5472
rect 5769 5408 5785 5472
rect 5849 5408 5865 5472
rect 5929 5408 5945 5472
rect 6009 5408 6017 5472
rect 5697 4966 6017 5408
rect 5697 4730 5739 4966
rect 5975 4730 6017 4966
rect 5697 4384 6017 4730
rect 5697 4320 5705 4384
rect 5769 4320 5785 4384
rect 5849 4320 5865 4384
rect 5929 4320 5945 4384
rect 6009 4320 6017 4384
rect 5697 3296 6017 4320
rect 5697 3232 5705 3296
rect 5769 3232 5785 3296
rect 5849 3232 5865 3296
rect 5929 3232 5945 3296
rect 6009 3232 6017 3296
rect 5697 3152 6017 3232
rect 5697 2916 5739 3152
rect 5975 2916 6017 3152
rect 5697 2208 6017 2916
rect 5697 2144 5705 2208
rect 5769 2144 5785 2208
rect 5849 2144 5865 2208
rect 5929 2144 5945 2208
rect 6009 2144 6017 2208
rect 5697 2128 6017 2144
<< via4 >>
rect 1936 6560 2172 6779
rect 1936 6543 1966 6560
rect 1966 6543 1982 6560
rect 1982 6543 2046 6560
rect 2046 6543 2062 6560
rect 2062 6543 2126 6560
rect 2126 6543 2142 6560
rect 2142 6543 2172 6560
rect 1936 4730 2172 4966
rect 1936 2916 2172 3152
rect 2887 5636 3123 5872
rect 2887 3840 3123 4059
rect 2887 3823 2917 3840
rect 2917 3823 2933 3840
rect 2933 3823 2997 3840
rect 2997 3823 3013 3840
rect 3013 3823 3077 3840
rect 3077 3823 3093 3840
rect 3093 3823 3123 3840
rect 3838 6560 4074 6779
rect 3838 6543 3868 6560
rect 3868 6543 3884 6560
rect 3884 6543 3948 6560
rect 3948 6543 3964 6560
rect 3964 6543 4028 6560
rect 4028 6543 4044 6560
rect 4044 6543 4074 6560
rect 3838 4730 4074 4966
rect 3838 2916 4074 3152
rect 4788 5636 5024 5872
rect 4788 3840 5024 4059
rect 4788 3823 4818 3840
rect 4818 3823 4834 3840
rect 4834 3823 4898 3840
rect 4898 3823 4914 3840
rect 4914 3823 4978 3840
rect 4978 3823 4994 3840
rect 4994 3823 5024 3840
rect 5739 6560 5975 6779
rect 5739 6543 5769 6560
rect 5769 6543 5785 6560
rect 5785 6543 5849 6560
rect 5849 6543 5865 6560
rect 5865 6543 5929 6560
rect 5929 6543 5945 6560
rect 5945 6543 5975 6560
rect 5739 4730 5975 4966
rect 5739 2916 5975 3152
<< metal5 >>
rect 1104 6779 6808 6821
rect 1104 6543 1936 6779
rect 2172 6543 3838 6779
rect 4074 6543 5739 6779
rect 5975 6543 6808 6779
rect 1104 6501 6808 6543
rect 1104 5872 6808 5915
rect 1104 5636 2887 5872
rect 3123 5636 4788 5872
rect 5024 5636 6808 5872
rect 1104 5594 6808 5636
rect 1104 4966 6808 5008
rect 1104 4730 1936 4966
rect 2172 4730 3838 4966
rect 4074 4730 5739 4966
rect 5975 4730 6808 4966
rect 1104 4688 6808 4730
rect 1104 4059 6808 4101
rect 1104 3823 2887 4059
rect 3123 3823 4788 4059
rect 5024 3823 6808 4059
rect 1104 3781 6808 3823
rect 1104 3152 6808 3195
rect 1104 2916 1936 3152
rect 2172 2916 3838 3152
rect 4074 2916 5739 3152
rect 5975 2916 6808 3152
rect 1104 2874 6808 2916
use sky130_fd_sc_hd__decap_4  FILLER_1_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 1932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8
timestamp 1623249630
transform 1 0 1840 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 1472 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform -1 0 1932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1623249630
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1623249630
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1623249630
transform 1 0 2576 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _25_
timestamp 1623249630
transform 1 0 2208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _19_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 2944 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 2300 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_1  _30_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 4232 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _31_
timestamp 1623249630
transform 1 0 4232 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25
timestamp 1623249630
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30
timestamp 1623249630
transform 1 0 3864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_29
timestamp 1623249630
transform 1 0 3772 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_33
timestamp 1623249630
transform 1 0 4140 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_42
timestamp 1623249630
transform 1 0 4968 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42
timestamp 1623249630
transform 1 0 4968 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _32_
timestamp 1623249630
transform 1 0 5336 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _28_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform -1 0 5796 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58
timestamp 1623249630
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54
timestamp 1623249630
transform 1 0 6072 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_22
timestamp 1623249630
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_21
timestamp 1623249630
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1623249630
transform -1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1623249630
transform -1 0 6808 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1623249630
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1623249630
transform -1 0 2024 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1623249630
transform 1 0 2392 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1623249630
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1623249630
transform 1 0 2024 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1623249630
transform 1 0 2668 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _27_
timestamp 1623249630
transform 1 0 3036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_23
timestamp 1623249630
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_25
timestamp 1623249630
transform 1 0 3404 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 3864 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_38
timestamp 1623249630
transform 1 0 4600 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1623249630
transform -1 0 6808 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1623249630
transform 1 0 5888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1623249630
transform 1 0 5520 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1623249630
transform 1 0 6164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform -1 0 3588 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1623249630
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1623249630
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 1623249630
transform 1 0 1380 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1623249630
transform 1 0 2392 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _35_
timestamp 1623249630
transform 1 0 3956 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1623249630
transform 1 0 3588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_40
timestamp 1623249630
transform 1 0 4784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _36_
timestamp 1623249630
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1623249630
transform -1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_24
timestamp 1623249630
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_53
timestamp 1623249630
transform 1 0 5980 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1623249630
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1623249630
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_15
timestamp 1623249630
transform 1 0 2484 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 3128 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _22_
timestamp 1623249630
transform -1 0 5060 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_25
timestamp 1623249630
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_21
timestamp 1623249630
transform 1 0 3036 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_25
timestamp 1623249630
transform 1 0 3404 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_30
timestamp 1623249630
transform 1 0 3864 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _29_
timestamp 1623249630
transform 1 0 5428 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1623249630
transform -1 0 6808 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_43
timestamp 1623249630
transform 1 0 5060 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_55
timestamp 1623249630
transform 1 0 6164 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _40_
timestamp 1623249630
transform -1 0 2852 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1623249630
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_19
timestamp 1623249630
transform 1 0 2852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 3404 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _26_
timestamp 1623249630
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1623249630
transform -1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_26
timestamp 1623249630
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_45
timestamp 1623249630
transform 1 0 5244 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_49
timestamp 1623249630
transform 1 0 5612 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_53
timestamp 1623249630
transform 1 0 5980 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1623249630
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1623249630
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1623249630
transform -1 0 2116 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1623249630
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1623249630
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_18
timestamp 1623249630
transform 1 0 2760 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_11
timestamp 1623249630
transform 1 0 2116 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_15
timestamp 1623249630
transform 1 0 2484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1623249630
transform -1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _23_
timestamp 1623249630
transform 1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1623249630
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__o221a_1  _24_
timestamp 1623249630
transform -1 0 5060 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _38_
timestamp 1623249630
transform -1 0 4600 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_27
timestamp 1623249630
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_25
timestamp 1623249630
transform 1 0 3404 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_30
timestamp 1623249630
transform 1 0 3864 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_38
timestamp 1623249630
transform 1 0 4600 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_51
timestamp 1623249630
transform 1 0 5796 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_50
timestamp 1623249630
transform 1 0 5704 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_43
timestamp 1623249630
transform 1 0 5060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _34_
timestamp 1623249630
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1623249630
transform 1 0 5428 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1623249630
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_58
timestamp 1623249630
transform 1 0 6440 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_28
timestamp 1623249630
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1623249630
transform -1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1623249630
transform -1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1623249630
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1623249630
transform -1 0 2760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1623249630
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1623249630
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _39_
timestamp 1623249630
transform 1 0 4232 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_29
timestamp 1623249630
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1623249630
transform -1 0 3404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_25
timestamp 1623249630
transform 1 0 3404 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_30
timestamp 1623249630
transform 1 0 3864 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1623249630
transform -1 0 6808 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_50
timestamp 1623249630
transform 1 0 5704 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1623249630
transform 1 0 6440 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1623249630
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1623249630
transform -1 0 2116 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output12
timestamp 1623249630
transform -1 0 2852 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1623249630
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_11
timestamp 1623249630
transform 1 0 2116 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_19
timestamp 1623249630
transform 1 0 2852 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_30
timestamp 1623249630
transform 1 0 3772 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1623249630
transform -1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1623249630
transform 1 0 3588 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_30
timestamp 1623249630
transform 1 0 3864 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_37
timestamp 1623249630
transform 1 0 4508 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1623249630
transform -1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_31
timestamp 1623249630
transform 1 0 6440 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1623249630
transform 1 0 5796 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1623249630
transform -1 0 5428 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp 1623249630
transform 1 0 5060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_47
timestamp 1623249630
transform 1 0 5428 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_54
timestamp 1623249630
transform 1 0 6072 0 1 7072
box -38 -48 406 592
<< labels >>
rlabel metal2 s 2318 0 2374 800 6 clk
port 0 nsew signal input
rlabel metal3 s 7199 6128 7999 6248 6 left
port 1 nsew signal input
rlabel metal2 s 7378 9343 7434 10143 6 parallelin[0]
port 2 nsew signal input
rlabel metal2 s 478 0 534 800 6 parallelin[1]
port 3 nsew signal input
rlabel metal3 s 7199 3408 7999 3528 6 parallelin[2]
port 4 nsew signal input
rlabel metal2 s 3698 9343 3754 10143 6 parallelin[3]
port 5 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 parallelout[0]
port 6 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 parallelout[1]
port 7 nsew signal tristate
rlabel metal2 s 1858 9343 1914 10143 6 parallelout[2]
port 8 nsew signal tristate
rlabel metal3 s 7199 688 7999 808 6 parallelout[3]
port 9 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 right
port 10 nsew signal input
rlabel metal2 s 5538 9343 5594 10143 6 rst
port 11 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 select[0]
port 12 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 select[1]
port 13 nsew signal input
rlabel metal4 s 5697 2128 6017 7664 6 VPWR
port 14 nsew power bidirectional
rlabel metal4 s 3796 2128 4116 7664 6 VPWR
port 15 nsew power bidirectional
rlabel metal4 s 1895 2128 2215 7664 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1104 6501 6808 6821 6 VPWR
port 17 nsew power bidirectional
rlabel metal5 s 1104 4688 6808 5008 6 VPWR
port 18 nsew power bidirectional
rlabel metal5 s 1104 2875 6808 3195 6 VPWR
port 19 nsew power bidirectional
rlabel metal4 s 4747 2128 5067 7664 6 VGND
port 20 nsew ground bidirectional
rlabel metal4 s 2845 2128 3165 7664 6 VGND
port 21 nsew ground bidirectional
rlabel metal5 s 1104 5595 6808 5915 6 VGND
port 22 nsew ground bidirectional
rlabel metal5 s 1104 3781 6808 4101 6 VGND
port 23 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 7999 10143
<< end >>
